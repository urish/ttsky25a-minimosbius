magic
tech sky130A
magscale 1 2
timestamp 1757105855
<< nwell >>
rect -358 -12269 358 12269
<< mvpmos >>
rect -100 7372 100 11972
rect -100 2536 100 7136
rect -100 -2300 100 2300
rect -100 -7136 100 -2536
rect -100 -11972 100 -7372
<< mvpdiff >>
rect -158 11960 -100 11972
rect -158 7384 -146 11960
rect -112 7384 -100 11960
rect -158 7372 -100 7384
rect 100 11960 158 11972
rect 100 7384 112 11960
rect 146 7384 158 11960
rect 100 7372 158 7384
rect -158 7124 -100 7136
rect -158 2548 -146 7124
rect -112 2548 -100 7124
rect -158 2536 -100 2548
rect 100 7124 158 7136
rect 100 2548 112 7124
rect 146 2548 158 7124
rect 100 2536 158 2548
rect -158 2288 -100 2300
rect -158 -2288 -146 2288
rect -112 -2288 -100 2288
rect -158 -2300 -100 -2288
rect 100 2288 158 2300
rect 100 -2288 112 2288
rect 146 -2288 158 2288
rect 100 -2300 158 -2288
rect -158 -2548 -100 -2536
rect -158 -7124 -146 -2548
rect -112 -7124 -100 -2548
rect -158 -7136 -100 -7124
rect 100 -2548 158 -2536
rect 100 -7124 112 -2548
rect 146 -7124 158 -2548
rect 100 -7136 158 -7124
rect -158 -7384 -100 -7372
rect -158 -11960 -146 -7384
rect -112 -11960 -100 -7384
rect -158 -11972 -100 -11960
rect 100 -7384 158 -7372
rect 100 -11960 112 -7384
rect 146 -11960 158 -7384
rect 100 -11972 158 -11960
<< mvpdiffc >>
rect -146 7384 -112 11960
rect 112 7384 146 11960
rect -146 2548 -112 7124
rect 112 2548 146 7124
rect -146 -2288 -112 2288
rect 112 -2288 146 2288
rect -146 -7124 -112 -2548
rect 112 -7124 146 -2548
rect -146 -11960 -112 -7384
rect 112 -11960 146 -7384
<< mvnsubdiff >>
rect -292 12191 292 12203
rect -292 12157 -184 12191
rect 184 12157 292 12191
rect -292 12145 292 12157
rect -292 12095 -234 12145
rect -292 -12095 -280 12095
rect -246 -12095 -234 12095
rect 234 12095 292 12145
rect -292 -12145 -234 -12095
rect 234 -12095 246 12095
rect 280 -12095 292 12095
rect 234 -12145 292 -12095
rect -292 -12157 292 -12145
rect -292 -12191 -184 -12157
rect 184 -12191 292 -12157
rect -292 -12203 292 -12191
<< mvnsubdiffcont >>
rect -184 12157 184 12191
rect -280 -12095 -246 12095
rect 246 -12095 280 12095
rect -184 -12191 184 -12157
<< poly >>
rect -100 12053 100 12069
rect -100 12019 -84 12053
rect 84 12019 100 12053
rect -100 11972 100 12019
rect -100 7325 100 7372
rect -100 7291 -84 7325
rect 84 7291 100 7325
rect -100 7275 100 7291
rect -100 7217 100 7233
rect -100 7183 -84 7217
rect 84 7183 100 7217
rect -100 7136 100 7183
rect -100 2489 100 2536
rect -100 2455 -84 2489
rect 84 2455 100 2489
rect -100 2439 100 2455
rect -100 2381 100 2397
rect -100 2347 -84 2381
rect 84 2347 100 2381
rect -100 2300 100 2347
rect -100 -2347 100 -2300
rect -100 -2381 -84 -2347
rect 84 -2381 100 -2347
rect -100 -2397 100 -2381
rect -100 -2455 100 -2439
rect -100 -2489 -84 -2455
rect 84 -2489 100 -2455
rect -100 -2536 100 -2489
rect -100 -7183 100 -7136
rect -100 -7217 -84 -7183
rect 84 -7217 100 -7183
rect -100 -7233 100 -7217
rect -100 -7291 100 -7275
rect -100 -7325 -84 -7291
rect 84 -7325 100 -7291
rect -100 -7372 100 -7325
rect -100 -12019 100 -11972
rect -100 -12053 -84 -12019
rect 84 -12053 100 -12019
rect -100 -12069 100 -12053
<< polycont >>
rect -84 12019 84 12053
rect -84 7291 84 7325
rect -84 7183 84 7217
rect -84 2455 84 2489
rect -84 2347 84 2381
rect -84 -2381 84 -2347
rect -84 -2489 84 -2455
rect -84 -7217 84 -7183
rect -84 -7325 84 -7291
rect -84 -12053 84 -12019
<< locali >>
rect -280 12157 -184 12191
rect 184 12157 280 12191
rect -280 12095 -246 12157
rect 246 12095 280 12157
rect -100 12019 -84 12053
rect 84 12019 100 12053
rect -146 11960 -112 11976
rect -146 7368 -112 7384
rect 112 11960 146 11976
rect 112 7368 146 7384
rect -100 7291 -84 7325
rect 84 7291 100 7325
rect -100 7183 -84 7217
rect 84 7183 100 7217
rect -146 7124 -112 7140
rect -146 2532 -112 2548
rect 112 7124 146 7140
rect 112 2532 146 2548
rect -100 2455 -84 2489
rect 84 2455 100 2489
rect -100 2347 -84 2381
rect 84 2347 100 2381
rect -146 2288 -112 2304
rect -146 -2304 -112 -2288
rect 112 2288 146 2304
rect 112 -2304 146 -2288
rect -100 -2381 -84 -2347
rect 84 -2381 100 -2347
rect -100 -2489 -84 -2455
rect 84 -2489 100 -2455
rect -146 -2548 -112 -2532
rect -146 -7140 -112 -7124
rect 112 -2548 146 -2532
rect 112 -7140 146 -7124
rect -100 -7217 -84 -7183
rect 84 -7217 100 -7183
rect -100 -7325 -84 -7291
rect 84 -7325 100 -7291
rect -146 -7384 -112 -7368
rect -146 -11976 -112 -11960
rect 112 -7384 146 -7368
rect 112 -11976 146 -11960
rect -100 -12053 -84 -12019
rect 84 -12053 100 -12019
rect -280 -12157 -246 -12095
rect 246 -12157 280 -12095
rect -280 -12191 -184 -12157
rect 184 -12191 280 -12157
<< viali >>
rect -84 12019 84 12053
rect -146 7384 -112 11960
rect 112 7384 146 11960
rect -84 7291 84 7325
rect -84 7183 84 7217
rect -146 2548 -112 7124
rect 112 2548 146 7124
rect -84 2455 84 2489
rect -84 2347 84 2381
rect -146 -2288 -112 2288
rect 112 -2288 146 2288
rect -84 -2381 84 -2347
rect -84 -2489 84 -2455
rect -146 -7124 -112 -2548
rect 112 -7124 146 -2548
rect -84 -7217 84 -7183
rect -84 -7325 84 -7291
rect -146 -11960 -112 -7384
rect 112 -11960 146 -7384
rect -84 -12053 84 -12019
<< metal1 >>
rect -96 12053 96 12059
rect -96 12019 -84 12053
rect 84 12019 96 12053
rect -96 12013 96 12019
rect -152 11960 -106 11972
rect -152 7384 -146 11960
rect -112 7384 -106 11960
rect -152 7372 -106 7384
rect 106 11960 152 11972
rect 106 7384 112 11960
rect 146 7384 152 11960
rect 106 7372 152 7384
rect -96 7325 96 7331
rect -96 7291 -84 7325
rect 84 7291 96 7325
rect -96 7285 96 7291
rect -96 7217 96 7223
rect -96 7183 -84 7217
rect 84 7183 96 7217
rect -96 7177 96 7183
rect -152 7124 -106 7136
rect -152 2548 -146 7124
rect -112 2548 -106 7124
rect -152 2536 -106 2548
rect 106 7124 152 7136
rect 106 2548 112 7124
rect 146 2548 152 7124
rect 106 2536 152 2548
rect -96 2489 96 2495
rect -96 2455 -84 2489
rect 84 2455 96 2489
rect -96 2449 96 2455
rect -96 2381 96 2387
rect -96 2347 -84 2381
rect 84 2347 96 2381
rect -96 2341 96 2347
rect -152 2288 -106 2300
rect -152 -2288 -146 2288
rect -112 -2288 -106 2288
rect -152 -2300 -106 -2288
rect 106 2288 152 2300
rect 106 -2288 112 2288
rect 146 -2288 152 2288
rect 106 -2300 152 -2288
rect -96 -2347 96 -2341
rect -96 -2381 -84 -2347
rect 84 -2381 96 -2347
rect -96 -2387 96 -2381
rect -96 -2455 96 -2449
rect -96 -2489 -84 -2455
rect 84 -2489 96 -2455
rect -96 -2495 96 -2489
rect -152 -2548 -106 -2536
rect -152 -7124 -146 -2548
rect -112 -7124 -106 -2548
rect -152 -7136 -106 -7124
rect 106 -2548 152 -2536
rect 106 -7124 112 -2548
rect 146 -7124 152 -2548
rect 106 -7136 152 -7124
rect -96 -7183 96 -7177
rect -96 -7217 -84 -7183
rect 84 -7217 96 -7183
rect -96 -7223 96 -7217
rect -96 -7291 96 -7285
rect -96 -7325 -84 -7291
rect 84 -7325 96 -7291
rect -96 -7331 96 -7325
rect -152 -7384 -106 -7372
rect -152 -11960 -146 -7384
rect -112 -11960 -106 -7384
rect -152 -11972 -106 -11960
rect 106 -7384 152 -7372
rect 106 -11960 112 -7384
rect 146 -11960 152 -7384
rect 106 -11972 152 -11960
rect -96 -12019 96 -12013
rect -96 -12053 -84 -12019
rect 84 -12053 96 -12019
rect -96 -12059 96 -12053
<< properties >>
string FIXED_BBOX -263 -12174 263 12174
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 23 l 1 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
