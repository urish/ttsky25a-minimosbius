magic
tech sky130A
magscale 1 2
timestamp 1757730208
<< pwell >>
rect -1621 -758 1621 758
<< mvnmos >>
rect -1393 -500 -1293 500
rect -1235 -500 -1135 500
rect -1077 -500 -977 500
rect -919 -500 -819 500
rect -761 -500 -661 500
rect -603 -500 -503 500
rect -445 -500 -345 500
rect -287 -500 -187 500
rect -129 -500 -29 500
rect 29 -500 129 500
rect 187 -500 287 500
rect 345 -500 445 500
rect 503 -500 603 500
rect 661 -500 761 500
rect 819 -500 919 500
rect 977 -500 1077 500
rect 1135 -500 1235 500
rect 1293 -500 1393 500
<< mvndiff >>
rect -1451 488 -1393 500
rect -1451 -488 -1439 488
rect -1405 -488 -1393 488
rect -1451 -500 -1393 -488
rect -1293 488 -1235 500
rect -1293 -488 -1281 488
rect -1247 -488 -1235 488
rect -1293 -500 -1235 -488
rect -1135 488 -1077 500
rect -1135 -488 -1123 488
rect -1089 -488 -1077 488
rect -1135 -500 -1077 -488
rect -977 488 -919 500
rect -977 -488 -965 488
rect -931 -488 -919 488
rect -977 -500 -919 -488
rect -819 488 -761 500
rect -819 -488 -807 488
rect -773 -488 -761 488
rect -819 -500 -761 -488
rect -661 488 -603 500
rect -661 -488 -649 488
rect -615 -488 -603 488
rect -661 -500 -603 -488
rect -503 488 -445 500
rect -503 -488 -491 488
rect -457 -488 -445 488
rect -503 -500 -445 -488
rect -345 488 -287 500
rect -345 -488 -333 488
rect -299 -488 -287 488
rect -345 -500 -287 -488
rect -187 488 -129 500
rect -187 -488 -175 488
rect -141 -488 -129 488
rect -187 -500 -129 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 129 488 187 500
rect 129 -488 141 488
rect 175 -488 187 488
rect 129 -500 187 -488
rect 287 488 345 500
rect 287 -488 299 488
rect 333 -488 345 488
rect 287 -500 345 -488
rect 445 488 503 500
rect 445 -488 457 488
rect 491 -488 503 488
rect 445 -500 503 -488
rect 603 488 661 500
rect 603 -488 615 488
rect 649 -488 661 488
rect 603 -500 661 -488
rect 761 488 819 500
rect 761 -488 773 488
rect 807 -488 819 488
rect 761 -500 819 -488
rect 919 488 977 500
rect 919 -488 931 488
rect 965 -488 977 488
rect 919 -500 977 -488
rect 1077 488 1135 500
rect 1077 -488 1089 488
rect 1123 -488 1135 488
rect 1077 -500 1135 -488
rect 1235 488 1293 500
rect 1235 -488 1247 488
rect 1281 -488 1293 488
rect 1235 -500 1293 -488
rect 1393 488 1451 500
rect 1393 -488 1405 488
rect 1439 -488 1451 488
rect 1393 -500 1451 -488
<< mvndiffc >>
rect -1439 -488 -1405 488
rect -1281 -488 -1247 488
rect -1123 -488 -1089 488
rect -965 -488 -931 488
rect -807 -488 -773 488
rect -649 -488 -615 488
rect -491 -488 -457 488
rect -333 -488 -299 488
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect 299 -488 333 488
rect 457 -488 491 488
rect 615 -488 649 488
rect 773 -488 807 488
rect 931 -488 965 488
rect 1089 -488 1123 488
rect 1247 -488 1281 488
rect 1405 -488 1439 488
<< mvpsubdiff >>
rect -1585 710 1585 722
rect -1585 676 -1477 710
rect 1477 676 1585 710
rect -1585 664 1585 676
rect -1585 614 -1527 664
rect -1585 -614 -1573 614
rect -1539 -614 -1527 614
rect 1527 614 1585 664
rect -1585 -664 -1527 -614
rect 1527 -614 1539 614
rect 1573 -614 1585 614
rect 1527 -664 1585 -614
rect -1585 -676 1585 -664
rect -1585 -710 -1477 -676
rect 1477 -710 1585 -676
rect -1585 -722 1585 -710
<< mvpsubdiffcont >>
rect -1477 676 1477 710
rect -1573 -614 -1539 614
rect 1539 -614 1573 614
rect -1477 -710 1477 -676
<< poly >>
rect -1393 572 -1293 588
rect -1393 538 -1377 572
rect -1309 538 -1293 572
rect -1393 500 -1293 538
rect -1235 572 -1135 588
rect -1235 538 -1219 572
rect -1151 538 -1135 572
rect -1235 500 -1135 538
rect -1077 572 -977 588
rect -1077 538 -1061 572
rect -993 538 -977 572
rect -1077 500 -977 538
rect -919 572 -819 588
rect -919 538 -903 572
rect -835 538 -819 572
rect -919 500 -819 538
rect -761 572 -661 588
rect -761 538 -745 572
rect -677 538 -661 572
rect -761 500 -661 538
rect -603 572 -503 588
rect -603 538 -587 572
rect -519 538 -503 572
rect -603 500 -503 538
rect -445 572 -345 588
rect -445 538 -429 572
rect -361 538 -345 572
rect -445 500 -345 538
rect -287 572 -187 588
rect -287 538 -271 572
rect -203 538 -187 572
rect -287 500 -187 538
rect -129 572 -29 588
rect -129 538 -113 572
rect -45 538 -29 572
rect -129 500 -29 538
rect 29 572 129 588
rect 29 538 45 572
rect 113 538 129 572
rect 29 500 129 538
rect 187 572 287 588
rect 187 538 203 572
rect 271 538 287 572
rect 187 500 287 538
rect 345 572 445 588
rect 345 538 361 572
rect 429 538 445 572
rect 345 500 445 538
rect 503 572 603 588
rect 503 538 519 572
rect 587 538 603 572
rect 503 500 603 538
rect 661 572 761 588
rect 661 538 677 572
rect 745 538 761 572
rect 661 500 761 538
rect 819 572 919 588
rect 819 538 835 572
rect 903 538 919 572
rect 819 500 919 538
rect 977 572 1077 588
rect 977 538 993 572
rect 1061 538 1077 572
rect 977 500 1077 538
rect 1135 572 1235 588
rect 1135 538 1151 572
rect 1219 538 1235 572
rect 1135 500 1235 538
rect 1293 572 1393 588
rect 1293 538 1309 572
rect 1377 538 1393 572
rect 1293 500 1393 538
rect -1393 -538 -1293 -500
rect -1393 -572 -1377 -538
rect -1309 -572 -1293 -538
rect -1393 -588 -1293 -572
rect -1235 -538 -1135 -500
rect -1235 -572 -1219 -538
rect -1151 -572 -1135 -538
rect -1235 -588 -1135 -572
rect -1077 -538 -977 -500
rect -1077 -572 -1061 -538
rect -993 -572 -977 -538
rect -1077 -588 -977 -572
rect -919 -538 -819 -500
rect -919 -572 -903 -538
rect -835 -572 -819 -538
rect -919 -588 -819 -572
rect -761 -538 -661 -500
rect -761 -572 -745 -538
rect -677 -572 -661 -538
rect -761 -588 -661 -572
rect -603 -538 -503 -500
rect -603 -572 -587 -538
rect -519 -572 -503 -538
rect -603 -588 -503 -572
rect -445 -538 -345 -500
rect -445 -572 -429 -538
rect -361 -572 -345 -538
rect -445 -588 -345 -572
rect -287 -538 -187 -500
rect -287 -572 -271 -538
rect -203 -572 -187 -538
rect -287 -588 -187 -572
rect -129 -538 -29 -500
rect -129 -572 -113 -538
rect -45 -572 -29 -538
rect -129 -588 -29 -572
rect 29 -538 129 -500
rect 29 -572 45 -538
rect 113 -572 129 -538
rect 29 -588 129 -572
rect 187 -538 287 -500
rect 187 -572 203 -538
rect 271 -572 287 -538
rect 187 -588 287 -572
rect 345 -538 445 -500
rect 345 -572 361 -538
rect 429 -572 445 -538
rect 345 -588 445 -572
rect 503 -538 603 -500
rect 503 -572 519 -538
rect 587 -572 603 -538
rect 503 -588 603 -572
rect 661 -538 761 -500
rect 661 -572 677 -538
rect 745 -572 761 -538
rect 661 -588 761 -572
rect 819 -538 919 -500
rect 819 -572 835 -538
rect 903 -572 919 -538
rect 819 -588 919 -572
rect 977 -538 1077 -500
rect 977 -572 993 -538
rect 1061 -572 1077 -538
rect 977 -588 1077 -572
rect 1135 -538 1235 -500
rect 1135 -572 1151 -538
rect 1219 -572 1235 -538
rect 1135 -588 1235 -572
rect 1293 -538 1393 -500
rect 1293 -572 1309 -538
rect 1377 -572 1393 -538
rect 1293 -588 1393 -572
<< polycont >>
rect -1377 538 -1309 572
rect -1219 538 -1151 572
rect -1061 538 -993 572
rect -903 538 -835 572
rect -745 538 -677 572
rect -587 538 -519 572
rect -429 538 -361 572
rect -271 538 -203 572
rect -113 538 -45 572
rect 45 538 113 572
rect 203 538 271 572
rect 361 538 429 572
rect 519 538 587 572
rect 677 538 745 572
rect 835 538 903 572
rect 993 538 1061 572
rect 1151 538 1219 572
rect 1309 538 1377 572
rect -1377 -572 -1309 -538
rect -1219 -572 -1151 -538
rect -1061 -572 -993 -538
rect -903 -572 -835 -538
rect -745 -572 -677 -538
rect -587 -572 -519 -538
rect -429 -572 -361 -538
rect -271 -572 -203 -538
rect -113 -572 -45 -538
rect 45 -572 113 -538
rect 203 -572 271 -538
rect 361 -572 429 -538
rect 519 -572 587 -538
rect 677 -572 745 -538
rect 835 -572 903 -538
rect 993 -572 1061 -538
rect 1151 -572 1219 -538
rect 1309 -572 1377 -538
<< locali >>
rect -1573 676 -1477 710
rect 1477 676 1573 710
rect -1573 614 -1539 676
rect 1539 614 1573 676
rect -1393 538 -1377 572
rect -1309 538 -1293 572
rect -1235 538 -1219 572
rect -1151 538 -1135 572
rect -1077 538 -1061 572
rect -993 538 -977 572
rect -919 538 -903 572
rect -835 538 -819 572
rect -761 538 -745 572
rect -677 538 -661 572
rect -603 538 -587 572
rect -519 538 -503 572
rect -445 538 -429 572
rect -361 538 -345 572
rect -287 538 -271 572
rect -203 538 -187 572
rect -129 538 -113 572
rect -45 538 -29 572
rect 29 538 45 572
rect 113 538 129 572
rect 187 538 203 572
rect 271 538 287 572
rect 345 538 361 572
rect 429 538 445 572
rect 503 538 519 572
rect 587 538 603 572
rect 661 538 677 572
rect 745 538 761 572
rect 819 538 835 572
rect 903 538 919 572
rect 977 538 993 572
rect 1061 538 1077 572
rect 1135 538 1151 572
rect 1219 538 1235 572
rect 1293 538 1309 572
rect 1377 538 1393 572
rect -1439 488 -1405 504
rect -1439 -504 -1405 -488
rect -1281 488 -1247 504
rect -1281 -504 -1247 -488
rect -1123 488 -1089 504
rect -1123 -504 -1089 -488
rect -965 488 -931 504
rect -965 -504 -931 -488
rect -807 488 -773 504
rect -807 -504 -773 -488
rect -649 488 -615 504
rect -649 -504 -615 -488
rect -491 488 -457 504
rect -491 -504 -457 -488
rect -333 488 -299 504
rect -333 -504 -299 -488
rect -175 488 -141 504
rect -175 -504 -141 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 141 488 175 504
rect 141 -504 175 -488
rect 299 488 333 504
rect 299 -504 333 -488
rect 457 488 491 504
rect 457 -504 491 -488
rect 615 488 649 504
rect 615 -504 649 -488
rect 773 488 807 504
rect 773 -504 807 -488
rect 931 488 965 504
rect 931 -504 965 -488
rect 1089 488 1123 504
rect 1089 -504 1123 -488
rect 1247 488 1281 504
rect 1247 -504 1281 -488
rect 1405 488 1439 504
rect 1405 -504 1439 -488
rect -1393 -572 -1377 -538
rect -1309 -572 -1293 -538
rect -1235 -572 -1219 -538
rect -1151 -572 -1135 -538
rect -1077 -572 -1061 -538
rect -993 -572 -977 -538
rect -919 -572 -903 -538
rect -835 -572 -819 -538
rect -761 -572 -745 -538
rect -677 -572 -661 -538
rect -603 -572 -587 -538
rect -519 -572 -503 -538
rect -445 -572 -429 -538
rect -361 -572 -345 -538
rect -287 -572 -271 -538
rect -203 -572 -187 -538
rect -129 -572 -113 -538
rect -45 -572 -29 -538
rect 29 -572 45 -538
rect 113 -572 129 -538
rect 187 -572 203 -538
rect 271 -572 287 -538
rect 345 -572 361 -538
rect 429 -572 445 -538
rect 503 -572 519 -538
rect 587 -572 603 -538
rect 661 -572 677 -538
rect 745 -572 761 -538
rect 819 -572 835 -538
rect 903 -572 919 -538
rect 977 -572 993 -538
rect 1061 -572 1077 -538
rect 1135 -572 1151 -538
rect 1219 -572 1235 -538
rect 1293 -572 1309 -538
rect 1377 -572 1393 -538
rect -1573 -676 -1539 -614
rect 1539 -676 1573 -614
rect -1573 -710 -1477 -676
rect 1477 -710 1573 -676
<< viali >>
rect -1377 538 -1309 572
rect -1219 538 -1151 572
rect -1061 538 -993 572
rect -903 538 -835 572
rect -745 538 -677 572
rect -587 538 -519 572
rect -429 538 -361 572
rect -271 538 -203 572
rect -113 538 -45 572
rect 45 538 113 572
rect 203 538 271 572
rect 361 538 429 572
rect 519 538 587 572
rect 677 538 745 572
rect 835 538 903 572
rect 993 538 1061 572
rect 1151 538 1219 572
rect 1309 538 1377 572
rect -1439 -488 -1405 488
rect -1281 -488 -1247 488
rect -1123 -488 -1089 488
rect -965 -488 -931 488
rect -807 -488 -773 488
rect -649 -488 -615 488
rect -491 -488 -457 488
rect -333 -488 -299 488
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect 299 -488 333 488
rect 457 -488 491 488
rect 615 -488 649 488
rect 773 -488 807 488
rect 931 -488 965 488
rect 1089 -488 1123 488
rect 1247 -488 1281 488
rect 1405 -488 1439 488
rect -1377 -572 -1309 -538
rect -1219 -572 -1151 -538
rect -1061 -572 -993 -538
rect -903 -572 -835 -538
rect -745 -572 -677 -538
rect -587 -572 -519 -538
rect -429 -572 -361 -538
rect -271 -572 -203 -538
rect -113 -572 -45 -538
rect 45 -572 113 -538
rect 203 -572 271 -538
rect 361 -572 429 -538
rect 519 -572 587 -538
rect 677 -572 745 -538
rect 835 -572 903 -538
rect 993 -572 1061 -538
rect 1151 -572 1219 -538
rect 1309 -572 1377 -538
<< metal1 >>
rect -1389 572 -1297 578
rect -1389 538 -1377 572
rect -1309 538 -1297 572
rect -1389 532 -1297 538
rect -1231 572 -1139 578
rect -1231 538 -1219 572
rect -1151 538 -1139 572
rect -1231 532 -1139 538
rect -1073 572 -981 578
rect -1073 538 -1061 572
rect -993 538 -981 572
rect -1073 532 -981 538
rect -915 572 -823 578
rect -915 538 -903 572
rect -835 538 -823 572
rect -915 532 -823 538
rect -757 572 -665 578
rect -757 538 -745 572
rect -677 538 -665 572
rect -757 532 -665 538
rect -599 572 -507 578
rect -599 538 -587 572
rect -519 538 -507 572
rect -599 532 -507 538
rect -441 572 -349 578
rect -441 538 -429 572
rect -361 538 -349 572
rect -441 532 -349 538
rect -283 572 -191 578
rect -283 538 -271 572
rect -203 538 -191 572
rect -283 532 -191 538
rect -125 572 -33 578
rect -125 538 -113 572
rect -45 538 -33 572
rect -125 532 -33 538
rect 33 572 125 578
rect 33 538 45 572
rect 113 538 125 572
rect 33 532 125 538
rect 191 572 283 578
rect 191 538 203 572
rect 271 538 283 572
rect 191 532 283 538
rect 349 572 441 578
rect 349 538 361 572
rect 429 538 441 572
rect 349 532 441 538
rect 507 572 599 578
rect 507 538 519 572
rect 587 538 599 572
rect 507 532 599 538
rect 665 572 757 578
rect 665 538 677 572
rect 745 538 757 572
rect 665 532 757 538
rect 823 572 915 578
rect 823 538 835 572
rect 903 538 915 572
rect 823 532 915 538
rect 981 572 1073 578
rect 981 538 993 572
rect 1061 538 1073 572
rect 981 532 1073 538
rect 1139 572 1231 578
rect 1139 538 1151 572
rect 1219 538 1231 572
rect 1139 532 1231 538
rect 1297 572 1389 578
rect 1297 538 1309 572
rect 1377 538 1389 572
rect 1297 532 1389 538
rect -1445 488 -1399 500
rect -1445 -488 -1439 488
rect -1405 -488 -1399 488
rect -1445 -500 -1399 -488
rect -1287 488 -1241 500
rect -1287 -488 -1281 488
rect -1247 -488 -1241 488
rect -1287 -500 -1241 -488
rect -1129 488 -1083 500
rect -1129 -488 -1123 488
rect -1089 -488 -1083 488
rect -1129 -500 -1083 -488
rect -971 488 -925 500
rect -971 -488 -965 488
rect -931 -488 -925 488
rect -971 -500 -925 -488
rect -813 488 -767 500
rect -813 -488 -807 488
rect -773 -488 -767 488
rect -813 -500 -767 -488
rect -655 488 -609 500
rect -655 -488 -649 488
rect -615 -488 -609 488
rect -655 -500 -609 -488
rect -497 488 -451 500
rect -497 -488 -491 488
rect -457 -488 -451 488
rect -497 -500 -451 -488
rect -339 488 -293 500
rect -339 -488 -333 488
rect -299 -488 -293 488
rect -339 -500 -293 -488
rect -181 488 -135 500
rect -181 -488 -175 488
rect -141 -488 -135 488
rect -181 -500 -135 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 135 488 181 500
rect 135 -488 141 488
rect 175 -488 181 488
rect 135 -500 181 -488
rect 293 488 339 500
rect 293 -488 299 488
rect 333 -488 339 488
rect 293 -500 339 -488
rect 451 488 497 500
rect 451 -488 457 488
rect 491 -488 497 488
rect 451 -500 497 -488
rect 609 488 655 500
rect 609 -488 615 488
rect 649 -488 655 488
rect 609 -500 655 -488
rect 767 488 813 500
rect 767 -488 773 488
rect 807 -488 813 488
rect 767 -500 813 -488
rect 925 488 971 500
rect 925 -488 931 488
rect 965 -488 971 488
rect 925 -500 971 -488
rect 1083 488 1129 500
rect 1083 -488 1089 488
rect 1123 -488 1129 488
rect 1083 -500 1129 -488
rect 1241 488 1287 500
rect 1241 -488 1247 488
rect 1281 -488 1287 488
rect 1241 -500 1287 -488
rect 1399 488 1445 500
rect 1399 -488 1405 488
rect 1439 -488 1445 488
rect 1399 -500 1445 -488
rect -1389 -538 -1297 -532
rect -1389 -572 -1377 -538
rect -1309 -572 -1297 -538
rect -1389 -578 -1297 -572
rect -1231 -538 -1139 -532
rect -1231 -572 -1219 -538
rect -1151 -572 -1139 -538
rect -1231 -578 -1139 -572
rect -1073 -538 -981 -532
rect -1073 -572 -1061 -538
rect -993 -572 -981 -538
rect -1073 -578 -981 -572
rect -915 -538 -823 -532
rect -915 -572 -903 -538
rect -835 -572 -823 -538
rect -915 -578 -823 -572
rect -757 -538 -665 -532
rect -757 -572 -745 -538
rect -677 -572 -665 -538
rect -757 -578 -665 -572
rect -599 -538 -507 -532
rect -599 -572 -587 -538
rect -519 -572 -507 -538
rect -599 -578 -507 -572
rect -441 -538 -349 -532
rect -441 -572 -429 -538
rect -361 -572 -349 -538
rect -441 -578 -349 -572
rect -283 -538 -191 -532
rect -283 -572 -271 -538
rect -203 -572 -191 -538
rect -283 -578 -191 -572
rect -125 -538 -33 -532
rect -125 -572 -113 -538
rect -45 -572 -33 -538
rect -125 -578 -33 -572
rect 33 -538 125 -532
rect 33 -572 45 -538
rect 113 -572 125 -538
rect 33 -578 125 -572
rect 191 -538 283 -532
rect 191 -572 203 -538
rect 271 -572 283 -538
rect 191 -578 283 -572
rect 349 -538 441 -532
rect 349 -572 361 -538
rect 429 -572 441 -538
rect 349 -578 441 -572
rect 507 -538 599 -532
rect 507 -572 519 -538
rect 587 -572 599 -538
rect 507 -578 599 -572
rect 665 -538 757 -532
rect 665 -572 677 -538
rect 745 -572 757 -538
rect 665 -578 757 -572
rect 823 -538 915 -532
rect 823 -572 835 -538
rect 903 -572 915 -538
rect 823 -578 915 -572
rect 981 -538 1073 -532
rect 981 -572 993 -538
rect 1061 -572 1073 -538
rect 981 -578 1073 -572
rect 1139 -538 1231 -532
rect 1139 -572 1151 -538
rect 1219 -572 1231 -538
rect 1139 -578 1231 -572
rect 1297 -538 1389 -532
rect 1297 -572 1309 -538
rect 1377 -572 1389 -538
rect 1297 -578 1389 -572
<< properties >>
string FIXED_BBOX -1556 -693 1556 693
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.50 m 1 nf 18 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
