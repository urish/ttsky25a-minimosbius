magic
tech sky130A
magscale 1 2
timestamp 1757730208
<< nwell >>
rect -3841 -2651 3841 2651
<< mvpmos >>
rect -3583 1354 -3383 2354
rect -3325 1354 -3125 2354
rect -3067 1354 -2867 2354
rect -2809 1354 -2609 2354
rect -2551 1354 -2351 2354
rect -2293 1354 -2093 2354
rect -2035 1354 -1835 2354
rect -1777 1354 -1577 2354
rect -1519 1354 -1319 2354
rect -1261 1354 -1061 2354
rect -1003 1354 -803 2354
rect -745 1354 -545 2354
rect -487 1354 -287 2354
rect -229 1354 -29 2354
rect 29 1354 229 2354
rect 287 1354 487 2354
rect 545 1354 745 2354
rect 803 1354 1003 2354
rect 1061 1354 1261 2354
rect 1319 1354 1519 2354
rect 1577 1354 1777 2354
rect 1835 1354 2035 2354
rect 2093 1354 2293 2354
rect 2351 1354 2551 2354
rect 2609 1354 2809 2354
rect 2867 1354 3067 2354
rect 3125 1354 3325 2354
rect 3383 1354 3583 2354
rect -3583 118 -3383 1118
rect -3325 118 -3125 1118
rect -3067 118 -2867 1118
rect -2809 118 -2609 1118
rect -2551 118 -2351 1118
rect -2293 118 -2093 1118
rect -2035 118 -1835 1118
rect -1777 118 -1577 1118
rect -1519 118 -1319 1118
rect -1261 118 -1061 1118
rect -1003 118 -803 1118
rect -745 118 -545 1118
rect -487 118 -287 1118
rect -229 118 -29 1118
rect 29 118 229 1118
rect 287 118 487 1118
rect 545 118 745 1118
rect 803 118 1003 1118
rect 1061 118 1261 1118
rect 1319 118 1519 1118
rect 1577 118 1777 1118
rect 1835 118 2035 1118
rect 2093 118 2293 1118
rect 2351 118 2551 1118
rect 2609 118 2809 1118
rect 2867 118 3067 1118
rect 3125 118 3325 1118
rect 3383 118 3583 1118
rect -3583 -1118 -3383 -118
rect -3325 -1118 -3125 -118
rect -3067 -1118 -2867 -118
rect -2809 -1118 -2609 -118
rect -2551 -1118 -2351 -118
rect -2293 -1118 -2093 -118
rect -2035 -1118 -1835 -118
rect -1777 -1118 -1577 -118
rect -1519 -1118 -1319 -118
rect -1261 -1118 -1061 -118
rect -1003 -1118 -803 -118
rect -745 -1118 -545 -118
rect -487 -1118 -287 -118
rect -229 -1118 -29 -118
rect 29 -1118 229 -118
rect 287 -1118 487 -118
rect 545 -1118 745 -118
rect 803 -1118 1003 -118
rect 1061 -1118 1261 -118
rect 1319 -1118 1519 -118
rect 1577 -1118 1777 -118
rect 1835 -1118 2035 -118
rect 2093 -1118 2293 -118
rect 2351 -1118 2551 -118
rect 2609 -1118 2809 -118
rect 2867 -1118 3067 -118
rect 3125 -1118 3325 -118
rect 3383 -1118 3583 -118
rect -3583 -2354 -3383 -1354
rect -3325 -2354 -3125 -1354
rect -3067 -2354 -2867 -1354
rect -2809 -2354 -2609 -1354
rect -2551 -2354 -2351 -1354
rect -2293 -2354 -2093 -1354
rect -2035 -2354 -1835 -1354
rect -1777 -2354 -1577 -1354
rect -1519 -2354 -1319 -1354
rect -1261 -2354 -1061 -1354
rect -1003 -2354 -803 -1354
rect -745 -2354 -545 -1354
rect -487 -2354 -287 -1354
rect -229 -2354 -29 -1354
rect 29 -2354 229 -1354
rect 287 -2354 487 -1354
rect 545 -2354 745 -1354
rect 803 -2354 1003 -1354
rect 1061 -2354 1261 -1354
rect 1319 -2354 1519 -1354
rect 1577 -2354 1777 -1354
rect 1835 -2354 2035 -1354
rect 2093 -2354 2293 -1354
rect 2351 -2354 2551 -1354
rect 2609 -2354 2809 -1354
rect 2867 -2354 3067 -1354
rect 3125 -2354 3325 -1354
rect 3383 -2354 3583 -1354
<< mvpdiff >>
rect -3641 2342 -3583 2354
rect -3641 1366 -3629 2342
rect -3595 1366 -3583 2342
rect -3641 1354 -3583 1366
rect -3383 2342 -3325 2354
rect -3383 1366 -3371 2342
rect -3337 1366 -3325 2342
rect -3383 1354 -3325 1366
rect -3125 2342 -3067 2354
rect -3125 1366 -3113 2342
rect -3079 1366 -3067 2342
rect -3125 1354 -3067 1366
rect -2867 2342 -2809 2354
rect -2867 1366 -2855 2342
rect -2821 1366 -2809 2342
rect -2867 1354 -2809 1366
rect -2609 2342 -2551 2354
rect -2609 1366 -2597 2342
rect -2563 1366 -2551 2342
rect -2609 1354 -2551 1366
rect -2351 2342 -2293 2354
rect -2351 1366 -2339 2342
rect -2305 1366 -2293 2342
rect -2351 1354 -2293 1366
rect -2093 2342 -2035 2354
rect -2093 1366 -2081 2342
rect -2047 1366 -2035 2342
rect -2093 1354 -2035 1366
rect -1835 2342 -1777 2354
rect -1835 1366 -1823 2342
rect -1789 1366 -1777 2342
rect -1835 1354 -1777 1366
rect -1577 2342 -1519 2354
rect -1577 1366 -1565 2342
rect -1531 1366 -1519 2342
rect -1577 1354 -1519 1366
rect -1319 2342 -1261 2354
rect -1319 1366 -1307 2342
rect -1273 1366 -1261 2342
rect -1319 1354 -1261 1366
rect -1061 2342 -1003 2354
rect -1061 1366 -1049 2342
rect -1015 1366 -1003 2342
rect -1061 1354 -1003 1366
rect -803 2342 -745 2354
rect -803 1366 -791 2342
rect -757 1366 -745 2342
rect -803 1354 -745 1366
rect -545 2342 -487 2354
rect -545 1366 -533 2342
rect -499 1366 -487 2342
rect -545 1354 -487 1366
rect -287 2342 -229 2354
rect -287 1366 -275 2342
rect -241 1366 -229 2342
rect -287 1354 -229 1366
rect -29 2342 29 2354
rect -29 1366 -17 2342
rect 17 1366 29 2342
rect -29 1354 29 1366
rect 229 2342 287 2354
rect 229 1366 241 2342
rect 275 1366 287 2342
rect 229 1354 287 1366
rect 487 2342 545 2354
rect 487 1366 499 2342
rect 533 1366 545 2342
rect 487 1354 545 1366
rect 745 2342 803 2354
rect 745 1366 757 2342
rect 791 1366 803 2342
rect 745 1354 803 1366
rect 1003 2342 1061 2354
rect 1003 1366 1015 2342
rect 1049 1366 1061 2342
rect 1003 1354 1061 1366
rect 1261 2342 1319 2354
rect 1261 1366 1273 2342
rect 1307 1366 1319 2342
rect 1261 1354 1319 1366
rect 1519 2342 1577 2354
rect 1519 1366 1531 2342
rect 1565 1366 1577 2342
rect 1519 1354 1577 1366
rect 1777 2342 1835 2354
rect 1777 1366 1789 2342
rect 1823 1366 1835 2342
rect 1777 1354 1835 1366
rect 2035 2342 2093 2354
rect 2035 1366 2047 2342
rect 2081 1366 2093 2342
rect 2035 1354 2093 1366
rect 2293 2342 2351 2354
rect 2293 1366 2305 2342
rect 2339 1366 2351 2342
rect 2293 1354 2351 1366
rect 2551 2342 2609 2354
rect 2551 1366 2563 2342
rect 2597 1366 2609 2342
rect 2551 1354 2609 1366
rect 2809 2342 2867 2354
rect 2809 1366 2821 2342
rect 2855 1366 2867 2342
rect 2809 1354 2867 1366
rect 3067 2342 3125 2354
rect 3067 1366 3079 2342
rect 3113 1366 3125 2342
rect 3067 1354 3125 1366
rect 3325 2342 3383 2354
rect 3325 1366 3337 2342
rect 3371 1366 3383 2342
rect 3325 1354 3383 1366
rect 3583 2342 3641 2354
rect 3583 1366 3595 2342
rect 3629 1366 3641 2342
rect 3583 1354 3641 1366
rect -3641 1106 -3583 1118
rect -3641 130 -3629 1106
rect -3595 130 -3583 1106
rect -3641 118 -3583 130
rect -3383 1106 -3325 1118
rect -3383 130 -3371 1106
rect -3337 130 -3325 1106
rect -3383 118 -3325 130
rect -3125 1106 -3067 1118
rect -3125 130 -3113 1106
rect -3079 130 -3067 1106
rect -3125 118 -3067 130
rect -2867 1106 -2809 1118
rect -2867 130 -2855 1106
rect -2821 130 -2809 1106
rect -2867 118 -2809 130
rect -2609 1106 -2551 1118
rect -2609 130 -2597 1106
rect -2563 130 -2551 1106
rect -2609 118 -2551 130
rect -2351 1106 -2293 1118
rect -2351 130 -2339 1106
rect -2305 130 -2293 1106
rect -2351 118 -2293 130
rect -2093 1106 -2035 1118
rect -2093 130 -2081 1106
rect -2047 130 -2035 1106
rect -2093 118 -2035 130
rect -1835 1106 -1777 1118
rect -1835 130 -1823 1106
rect -1789 130 -1777 1106
rect -1835 118 -1777 130
rect -1577 1106 -1519 1118
rect -1577 130 -1565 1106
rect -1531 130 -1519 1106
rect -1577 118 -1519 130
rect -1319 1106 -1261 1118
rect -1319 130 -1307 1106
rect -1273 130 -1261 1106
rect -1319 118 -1261 130
rect -1061 1106 -1003 1118
rect -1061 130 -1049 1106
rect -1015 130 -1003 1106
rect -1061 118 -1003 130
rect -803 1106 -745 1118
rect -803 130 -791 1106
rect -757 130 -745 1106
rect -803 118 -745 130
rect -545 1106 -487 1118
rect -545 130 -533 1106
rect -499 130 -487 1106
rect -545 118 -487 130
rect -287 1106 -229 1118
rect -287 130 -275 1106
rect -241 130 -229 1106
rect -287 118 -229 130
rect -29 1106 29 1118
rect -29 130 -17 1106
rect 17 130 29 1106
rect -29 118 29 130
rect 229 1106 287 1118
rect 229 130 241 1106
rect 275 130 287 1106
rect 229 118 287 130
rect 487 1106 545 1118
rect 487 130 499 1106
rect 533 130 545 1106
rect 487 118 545 130
rect 745 1106 803 1118
rect 745 130 757 1106
rect 791 130 803 1106
rect 745 118 803 130
rect 1003 1106 1061 1118
rect 1003 130 1015 1106
rect 1049 130 1061 1106
rect 1003 118 1061 130
rect 1261 1106 1319 1118
rect 1261 130 1273 1106
rect 1307 130 1319 1106
rect 1261 118 1319 130
rect 1519 1106 1577 1118
rect 1519 130 1531 1106
rect 1565 130 1577 1106
rect 1519 118 1577 130
rect 1777 1106 1835 1118
rect 1777 130 1789 1106
rect 1823 130 1835 1106
rect 1777 118 1835 130
rect 2035 1106 2093 1118
rect 2035 130 2047 1106
rect 2081 130 2093 1106
rect 2035 118 2093 130
rect 2293 1106 2351 1118
rect 2293 130 2305 1106
rect 2339 130 2351 1106
rect 2293 118 2351 130
rect 2551 1106 2609 1118
rect 2551 130 2563 1106
rect 2597 130 2609 1106
rect 2551 118 2609 130
rect 2809 1106 2867 1118
rect 2809 130 2821 1106
rect 2855 130 2867 1106
rect 2809 118 2867 130
rect 3067 1106 3125 1118
rect 3067 130 3079 1106
rect 3113 130 3125 1106
rect 3067 118 3125 130
rect 3325 1106 3383 1118
rect 3325 130 3337 1106
rect 3371 130 3383 1106
rect 3325 118 3383 130
rect 3583 1106 3641 1118
rect 3583 130 3595 1106
rect 3629 130 3641 1106
rect 3583 118 3641 130
rect -3641 -130 -3583 -118
rect -3641 -1106 -3629 -130
rect -3595 -1106 -3583 -130
rect -3641 -1118 -3583 -1106
rect -3383 -130 -3325 -118
rect -3383 -1106 -3371 -130
rect -3337 -1106 -3325 -130
rect -3383 -1118 -3325 -1106
rect -3125 -130 -3067 -118
rect -3125 -1106 -3113 -130
rect -3079 -1106 -3067 -130
rect -3125 -1118 -3067 -1106
rect -2867 -130 -2809 -118
rect -2867 -1106 -2855 -130
rect -2821 -1106 -2809 -130
rect -2867 -1118 -2809 -1106
rect -2609 -130 -2551 -118
rect -2609 -1106 -2597 -130
rect -2563 -1106 -2551 -130
rect -2609 -1118 -2551 -1106
rect -2351 -130 -2293 -118
rect -2351 -1106 -2339 -130
rect -2305 -1106 -2293 -130
rect -2351 -1118 -2293 -1106
rect -2093 -130 -2035 -118
rect -2093 -1106 -2081 -130
rect -2047 -1106 -2035 -130
rect -2093 -1118 -2035 -1106
rect -1835 -130 -1777 -118
rect -1835 -1106 -1823 -130
rect -1789 -1106 -1777 -130
rect -1835 -1118 -1777 -1106
rect -1577 -130 -1519 -118
rect -1577 -1106 -1565 -130
rect -1531 -1106 -1519 -130
rect -1577 -1118 -1519 -1106
rect -1319 -130 -1261 -118
rect -1319 -1106 -1307 -130
rect -1273 -1106 -1261 -130
rect -1319 -1118 -1261 -1106
rect -1061 -130 -1003 -118
rect -1061 -1106 -1049 -130
rect -1015 -1106 -1003 -130
rect -1061 -1118 -1003 -1106
rect -803 -130 -745 -118
rect -803 -1106 -791 -130
rect -757 -1106 -745 -130
rect -803 -1118 -745 -1106
rect -545 -130 -487 -118
rect -545 -1106 -533 -130
rect -499 -1106 -487 -130
rect -545 -1118 -487 -1106
rect -287 -130 -229 -118
rect -287 -1106 -275 -130
rect -241 -1106 -229 -130
rect -287 -1118 -229 -1106
rect -29 -130 29 -118
rect -29 -1106 -17 -130
rect 17 -1106 29 -130
rect -29 -1118 29 -1106
rect 229 -130 287 -118
rect 229 -1106 241 -130
rect 275 -1106 287 -130
rect 229 -1118 287 -1106
rect 487 -130 545 -118
rect 487 -1106 499 -130
rect 533 -1106 545 -130
rect 487 -1118 545 -1106
rect 745 -130 803 -118
rect 745 -1106 757 -130
rect 791 -1106 803 -130
rect 745 -1118 803 -1106
rect 1003 -130 1061 -118
rect 1003 -1106 1015 -130
rect 1049 -1106 1061 -130
rect 1003 -1118 1061 -1106
rect 1261 -130 1319 -118
rect 1261 -1106 1273 -130
rect 1307 -1106 1319 -130
rect 1261 -1118 1319 -1106
rect 1519 -130 1577 -118
rect 1519 -1106 1531 -130
rect 1565 -1106 1577 -130
rect 1519 -1118 1577 -1106
rect 1777 -130 1835 -118
rect 1777 -1106 1789 -130
rect 1823 -1106 1835 -130
rect 1777 -1118 1835 -1106
rect 2035 -130 2093 -118
rect 2035 -1106 2047 -130
rect 2081 -1106 2093 -130
rect 2035 -1118 2093 -1106
rect 2293 -130 2351 -118
rect 2293 -1106 2305 -130
rect 2339 -1106 2351 -130
rect 2293 -1118 2351 -1106
rect 2551 -130 2609 -118
rect 2551 -1106 2563 -130
rect 2597 -1106 2609 -130
rect 2551 -1118 2609 -1106
rect 2809 -130 2867 -118
rect 2809 -1106 2821 -130
rect 2855 -1106 2867 -130
rect 2809 -1118 2867 -1106
rect 3067 -130 3125 -118
rect 3067 -1106 3079 -130
rect 3113 -1106 3125 -130
rect 3067 -1118 3125 -1106
rect 3325 -130 3383 -118
rect 3325 -1106 3337 -130
rect 3371 -1106 3383 -130
rect 3325 -1118 3383 -1106
rect 3583 -130 3641 -118
rect 3583 -1106 3595 -130
rect 3629 -1106 3641 -130
rect 3583 -1118 3641 -1106
rect -3641 -1366 -3583 -1354
rect -3641 -2342 -3629 -1366
rect -3595 -2342 -3583 -1366
rect -3641 -2354 -3583 -2342
rect -3383 -1366 -3325 -1354
rect -3383 -2342 -3371 -1366
rect -3337 -2342 -3325 -1366
rect -3383 -2354 -3325 -2342
rect -3125 -1366 -3067 -1354
rect -3125 -2342 -3113 -1366
rect -3079 -2342 -3067 -1366
rect -3125 -2354 -3067 -2342
rect -2867 -1366 -2809 -1354
rect -2867 -2342 -2855 -1366
rect -2821 -2342 -2809 -1366
rect -2867 -2354 -2809 -2342
rect -2609 -1366 -2551 -1354
rect -2609 -2342 -2597 -1366
rect -2563 -2342 -2551 -1366
rect -2609 -2354 -2551 -2342
rect -2351 -1366 -2293 -1354
rect -2351 -2342 -2339 -1366
rect -2305 -2342 -2293 -1366
rect -2351 -2354 -2293 -2342
rect -2093 -1366 -2035 -1354
rect -2093 -2342 -2081 -1366
rect -2047 -2342 -2035 -1366
rect -2093 -2354 -2035 -2342
rect -1835 -1366 -1777 -1354
rect -1835 -2342 -1823 -1366
rect -1789 -2342 -1777 -1366
rect -1835 -2354 -1777 -2342
rect -1577 -1366 -1519 -1354
rect -1577 -2342 -1565 -1366
rect -1531 -2342 -1519 -1366
rect -1577 -2354 -1519 -2342
rect -1319 -1366 -1261 -1354
rect -1319 -2342 -1307 -1366
rect -1273 -2342 -1261 -1366
rect -1319 -2354 -1261 -2342
rect -1061 -1366 -1003 -1354
rect -1061 -2342 -1049 -1366
rect -1015 -2342 -1003 -1366
rect -1061 -2354 -1003 -2342
rect -803 -1366 -745 -1354
rect -803 -2342 -791 -1366
rect -757 -2342 -745 -1366
rect -803 -2354 -745 -2342
rect -545 -1366 -487 -1354
rect -545 -2342 -533 -1366
rect -499 -2342 -487 -1366
rect -545 -2354 -487 -2342
rect -287 -1366 -229 -1354
rect -287 -2342 -275 -1366
rect -241 -2342 -229 -1366
rect -287 -2354 -229 -2342
rect -29 -1366 29 -1354
rect -29 -2342 -17 -1366
rect 17 -2342 29 -1366
rect -29 -2354 29 -2342
rect 229 -1366 287 -1354
rect 229 -2342 241 -1366
rect 275 -2342 287 -1366
rect 229 -2354 287 -2342
rect 487 -1366 545 -1354
rect 487 -2342 499 -1366
rect 533 -2342 545 -1366
rect 487 -2354 545 -2342
rect 745 -1366 803 -1354
rect 745 -2342 757 -1366
rect 791 -2342 803 -1366
rect 745 -2354 803 -2342
rect 1003 -1366 1061 -1354
rect 1003 -2342 1015 -1366
rect 1049 -2342 1061 -1366
rect 1003 -2354 1061 -2342
rect 1261 -1366 1319 -1354
rect 1261 -2342 1273 -1366
rect 1307 -2342 1319 -1366
rect 1261 -2354 1319 -2342
rect 1519 -1366 1577 -1354
rect 1519 -2342 1531 -1366
rect 1565 -2342 1577 -1366
rect 1519 -2354 1577 -2342
rect 1777 -1366 1835 -1354
rect 1777 -2342 1789 -1366
rect 1823 -2342 1835 -1366
rect 1777 -2354 1835 -2342
rect 2035 -1366 2093 -1354
rect 2035 -2342 2047 -1366
rect 2081 -2342 2093 -1366
rect 2035 -2354 2093 -2342
rect 2293 -1366 2351 -1354
rect 2293 -2342 2305 -1366
rect 2339 -2342 2351 -1366
rect 2293 -2354 2351 -2342
rect 2551 -1366 2609 -1354
rect 2551 -2342 2563 -1366
rect 2597 -2342 2609 -1366
rect 2551 -2354 2609 -2342
rect 2809 -1366 2867 -1354
rect 2809 -2342 2821 -1366
rect 2855 -2342 2867 -1366
rect 2809 -2354 2867 -2342
rect 3067 -1366 3125 -1354
rect 3067 -2342 3079 -1366
rect 3113 -2342 3125 -1366
rect 3067 -2354 3125 -2342
rect 3325 -1366 3383 -1354
rect 3325 -2342 3337 -1366
rect 3371 -2342 3383 -1366
rect 3325 -2354 3383 -2342
rect 3583 -1366 3641 -1354
rect 3583 -2342 3595 -1366
rect 3629 -2342 3641 -1366
rect 3583 -2354 3641 -2342
<< mvpdiffc >>
rect -3629 1366 -3595 2342
rect -3371 1366 -3337 2342
rect -3113 1366 -3079 2342
rect -2855 1366 -2821 2342
rect -2597 1366 -2563 2342
rect -2339 1366 -2305 2342
rect -2081 1366 -2047 2342
rect -1823 1366 -1789 2342
rect -1565 1366 -1531 2342
rect -1307 1366 -1273 2342
rect -1049 1366 -1015 2342
rect -791 1366 -757 2342
rect -533 1366 -499 2342
rect -275 1366 -241 2342
rect -17 1366 17 2342
rect 241 1366 275 2342
rect 499 1366 533 2342
rect 757 1366 791 2342
rect 1015 1366 1049 2342
rect 1273 1366 1307 2342
rect 1531 1366 1565 2342
rect 1789 1366 1823 2342
rect 2047 1366 2081 2342
rect 2305 1366 2339 2342
rect 2563 1366 2597 2342
rect 2821 1366 2855 2342
rect 3079 1366 3113 2342
rect 3337 1366 3371 2342
rect 3595 1366 3629 2342
rect -3629 130 -3595 1106
rect -3371 130 -3337 1106
rect -3113 130 -3079 1106
rect -2855 130 -2821 1106
rect -2597 130 -2563 1106
rect -2339 130 -2305 1106
rect -2081 130 -2047 1106
rect -1823 130 -1789 1106
rect -1565 130 -1531 1106
rect -1307 130 -1273 1106
rect -1049 130 -1015 1106
rect -791 130 -757 1106
rect -533 130 -499 1106
rect -275 130 -241 1106
rect -17 130 17 1106
rect 241 130 275 1106
rect 499 130 533 1106
rect 757 130 791 1106
rect 1015 130 1049 1106
rect 1273 130 1307 1106
rect 1531 130 1565 1106
rect 1789 130 1823 1106
rect 2047 130 2081 1106
rect 2305 130 2339 1106
rect 2563 130 2597 1106
rect 2821 130 2855 1106
rect 3079 130 3113 1106
rect 3337 130 3371 1106
rect 3595 130 3629 1106
rect -3629 -1106 -3595 -130
rect -3371 -1106 -3337 -130
rect -3113 -1106 -3079 -130
rect -2855 -1106 -2821 -130
rect -2597 -1106 -2563 -130
rect -2339 -1106 -2305 -130
rect -2081 -1106 -2047 -130
rect -1823 -1106 -1789 -130
rect -1565 -1106 -1531 -130
rect -1307 -1106 -1273 -130
rect -1049 -1106 -1015 -130
rect -791 -1106 -757 -130
rect -533 -1106 -499 -130
rect -275 -1106 -241 -130
rect -17 -1106 17 -130
rect 241 -1106 275 -130
rect 499 -1106 533 -130
rect 757 -1106 791 -130
rect 1015 -1106 1049 -130
rect 1273 -1106 1307 -130
rect 1531 -1106 1565 -130
rect 1789 -1106 1823 -130
rect 2047 -1106 2081 -130
rect 2305 -1106 2339 -130
rect 2563 -1106 2597 -130
rect 2821 -1106 2855 -130
rect 3079 -1106 3113 -130
rect 3337 -1106 3371 -130
rect 3595 -1106 3629 -130
rect -3629 -2342 -3595 -1366
rect -3371 -2342 -3337 -1366
rect -3113 -2342 -3079 -1366
rect -2855 -2342 -2821 -1366
rect -2597 -2342 -2563 -1366
rect -2339 -2342 -2305 -1366
rect -2081 -2342 -2047 -1366
rect -1823 -2342 -1789 -1366
rect -1565 -2342 -1531 -1366
rect -1307 -2342 -1273 -1366
rect -1049 -2342 -1015 -1366
rect -791 -2342 -757 -1366
rect -533 -2342 -499 -1366
rect -275 -2342 -241 -1366
rect -17 -2342 17 -1366
rect 241 -2342 275 -1366
rect 499 -2342 533 -1366
rect 757 -2342 791 -1366
rect 1015 -2342 1049 -1366
rect 1273 -2342 1307 -1366
rect 1531 -2342 1565 -1366
rect 1789 -2342 1823 -1366
rect 2047 -2342 2081 -1366
rect 2305 -2342 2339 -1366
rect 2563 -2342 2597 -1366
rect 2821 -2342 2855 -1366
rect 3079 -2342 3113 -1366
rect 3337 -2342 3371 -1366
rect 3595 -2342 3629 -1366
<< mvnsubdiff >>
rect -3775 2573 3775 2585
rect -3775 2539 -3667 2573
rect 3667 2539 3775 2573
rect -3775 2527 3775 2539
rect -3775 2477 -3717 2527
rect -3775 -2477 -3763 2477
rect -3729 -2477 -3717 2477
rect 3717 2477 3775 2527
rect -3775 -2527 -3717 -2477
rect 3717 -2477 3729 2477
rect 3763 -2477 3775 2477
rect 3717 -2527 3775 -2477
rect -3775 -2539 3775 -2527
rect -3775 -2573 -3667 -2539
rect 3667 -2573 3775 -2539
rect -3775 -2585 3775 -2573
<< mvnsubdiffcont >>
rect -3667 2539 3667 2573
rect -3763 -2477 -3729 2477
rect 3729 -2477 3763 2477
rect -3667 -2573 3667 -2539
<< poly >>
rect -3583 2435 -3383 2451
rect -3583 2401 -3567 2435
rect -3399 2401 -3383 2435
rect -3583 2354 -3383 2401
rect -3325 2435 -3125 2451
rect -3325 2401 -3309 2435
rect -3141 2401 -3125 2435
rect -3325 2354 -3125 2401
rect -3067 2435 -2867 2451
rect -3067 2401 -3051 2435
rect -2883 2401 -2867 2435
rect -3067 2354 -2867 2401
rect -2809 2435 -2609 2451
rect -2809 2401 -2793 2435
rect -2625 2401 -2609 2435
rect -2809 2354 -2609 2401
rect -2551 2435 -2351 2451
rect -2551 2401 -2535 2435
rect -2367 2401 -2351 2435
rect -2551 2354 -2351 2401
rect -2293 2435 -2093 2451
rect -2293 2401 -2277 2435
rect -2109 2401 -2093 2435
rect -2293 2354 -2093 2401
rect -2035 2435 -1835 2451
rect -2035 2401 -2019 2435
rect -1851 2401 -1835 2435
rect -2035 2354 -1835 2401
rect -1777 2435 -1577 2451
rect -1777 2401 -1761 2435
rect -1593 2401 -1577 2435
rect -1777 2354 -1577 2401
rect -1519 2435 -1319 2451
rect -1519 2401 -1503 2435
rect -1335 2401 -1319 2435
rect -1519 2354 -1319 2401
rect -1261 2435 -1061 2451
rect -1261 2401 -1245 2435
rect -1077 2401 -1061 2435
rect -1261 2354 -1061 2401
rect -1003 2435 -803 2451
rect -1003 2401 -987 2435
rect -819 2401 -803 2435
rect -1003 2354 -803 2401
rect -745 2435 -545 2451
rect -745 2401 -729 2435
rect -561 2401 -545 2435
rect -745 2354 -545 2401
rect -487 2435 -287 2451
rect -487 2401 -471 2435
rect -303 2401 -287 2435
rect -487 2354 -287 2401
rect -229 2435 -29 2451
rect -229 2401 -213 2435
rect -45 2401 -29 2435
rect -229 2354 -29 2401
rect 29 2435 229 2451
rect 29 2401 45 2435
rect 213 2401 229 2435
rect 29 2354 229 2401
rect 287 2435 487 2451
rect 287 2401 303 2435
rect 471 2401 487 2435
rect 287 2354 487 2401
rect 545 2435 745 2451
rect 545 2401 561 2435
rect 729 2401 745 2435
rect 545 2354 745 2401
rect 803 2435 1003 2451
rect 803 2401 819 2435
rect 987 2401 1003 2435
rect 803 2354 1003 2401
rect 1061 2435 1261 2451
rect 1061 2401 1077 2435
rect 1245 2401 1261 2435
rect 1061 2354 1261 2401
rect 1319 2435 1519 2451
rect 1319 2401 1335 2435
rect 1503 2401 1519 2435
rect 1319 2354 1519 2401
rect 1577 2435 1777 2451
rect 1577 2401 1593 2435
rect 1761 2401 1777 2435
rect 1577 2354 1777 2401
rect 1835 2435 2035 2451
rect 1835 2401 1851 2435
rect 2019 2401 2035 2435
rect 1835 2354 2035 2401
rect 2093 2435 2293 2451
rect 2093 2401 2109 2435
rect 2277 2401 2293 2435
rect 2093 2354 2293 2401
rect 2351 2435 2551 2451
rect 2351 2401 2367 2435
rect 2535 2401 2551 2435
rect 2351 2354 2551 2401
rect 2609 2435 2809 2451
rect 2609 2401 2625 2435
rect 2793 2401 2809 2435
rect 2609 2354 2809 2401
rect 2867 2435 3067 2451
rect 2867 2401 2883 2435
rect 3051 2401 3067 2435
rect 2867 2354 3067 2401
rect 3125 2435 3325 2451
rect 3125 2401 3141 2435
rect 3309 2401 3325 2435
rect 3125 2354 3325 2401
rect 3383 2435 3583 2451
rect 3383 2401 3399 2435
rect 3567 2401 3583 2435
rect 3383 2354 3583 2401
rect -3583 1307 -3383 1354
rect -3583 1273 -3567 1307
rect -3399 1273 -3383 1307
rect -3583 1257 -3383 1273
rect -3325 1307 -3125 1354
rect -3325 1273 -3309 1307
rect -3141 1273 -3125 1307
rect -3325 1257 -3125 1273
rect -3067 1307 -2867 1354
rect -3067 1273 -3051 1307
rect -2883 1273 -2867 1307
rect -3067 1257 -2867 1273
rect -2809 1307 -2609 1354
rect -2809 1273 -2793 1307
rect -2625 1273 -2609 1307
rect -2809 1257 -2609 1273
rect -2551 1307 -2351 1354
rect -2551 1273 -2535 1307
rect -2367 1273 -2351 1307
rect -2551 1257 -2351 1273
rect -2293 1307 -2093 1354
rect -2293 1273 -2277 1307
rect -2109 1273 -2093 1307
rect -2293 1257 -2093 1273
rect -2035 1307 -1835 1354
rect -2035 1273 -2019 1307
rect -1851 1273 -1835 1307
rect -2035 1257 -1835 1273
rect -1777 1307 -1577 1354
rect -1777 1273 -1761 1307
rect -1593 1273 -1577 1307
rect -1777 1257 -1577 1273
rect -1519 1307 -1319 1354
rect -1519 1273 -1503 1307
rect -1335 1273 -1319 1307
rect -1519 1257 -1319 1273
rect -1261 1307 -1061 1354
rect -1261 1273 -1245 1307
rect -1077 1273 -1061 1307
rect -1261 1257 -1061 1273
rect -1003 1307 -803 1354
rect -1003 1273 -987 1307
rect -819 1273 -803 1307
rect -1003 1257 -803 1273
rect -745 1307 -545 1354
rect -745 1273 -729 1307
rect -561 1273 -545 1307
rect -745 1257 -545 1273
rect -487 1307 -287 1354
rect -487 1273 -471 1307
rect -303 1273 -287 1307
rect -487 1257 -287 1273
rect -229 1307 -29 1354
rect -229 1273 -213 1307
rect -45 1273 -29 1307
rect -229 1257 -29 1273
rect 29 1307 229 1354
rect 29 1273 45 1307
rect 213 1273 229 1307
rect 29 1257 229 1273
rect 287 1307 487 1354
rect 287 1273 303 1307
rect 471 1273 487 1307
rect 287 1257 487 1273
rect 545 1307 745 1354
rect 545 1273 561 1307
rect 729 1273 745 1307
rect 545 1257 745 1273
rect 803 1307 1003 1354
rect 803 1273 819 1307
rect 987 1273 1003 1307
rect 803 1257 1003 1273
rect 1061 1307 1261 1354
rect 1061 1273 1077 1307
rect 1245 1273 1261 1307
rect 1061 1257 1261 1273
rect 1319 1307 1519 1354
rect 1319 1273 1335 1307
rect 1503 1273 1519 1307
rect 1319 1257 1519 1273
rect 1577 1307 1777 1354
rect 1577 1273 1593 1307
rect 1761 1273 1777 1307
rect 1577 1257 1777 1273
rect 1835 1307 2035 1354
rect 1835 1273 1851 1307
rect 2019 1273 2035 1307
rect 1835 1257 2035 1273
rect 2093 1307 2293 1354
rect 2093 1273 2109 1307
rect 2277 1273 2293 1307
rect 2093 1257 2293 1273
rect 2351 1307 2551 1354
rect 2351 1273 2367 1307
rect 2535 1273 2551 1307
rect 2351 1257 2551 1273
rect 2609 1307 2809 1354
rect 2609 1273 2625 1307
rect 2793 1273 2809 1307
rect 2609 1257 2809 1273
rect 2867 1307 3067 1354
rect 2867 1273 2883 1307
rect 3051 1273 3067 1307
rect 2867 1257 3067 1273
rect 3125 1307 3325 1354
rect 3125 1273 3141 1307
rect 3309 1273 3325 1307
rect 3125 1257 3325 1273
rect 3383 1307 3583 1354
rect 3383 1273 3399 1307
rect 3567 1273 3583 1307
rect 3383 1257 3583 1273
rect -3583 1199 -3383 1215
rect -3583 1165 -3567 1199
rect -3399 1165 -3383 1199
rect -3583 1118 -3383 1165
rect -3325 1199 -3125 1215
rect -3325 1165 -3309 1199
rect -3141 1165 -3125 1199
rect -3325 1118 -3125 1165
rect -3067 1199 -2867 1215
rect -3067 1165 -3051 1199
rect -2883 1165 -2867 1199
rect -3067 1118 -2867 1165
rect -2809 1199 -2609 1215
rect -2809 1165 -2793 1199
rect -2625 1165 -2609 1199
rect -2809 1118 -2609 1165
rect -2551 1199 -2351 1215
rect -2551 1165 -2535 1199
rect -2367 1165 -2351 1199
rect -2551 1118 -2351 1165
rect -2293 1199 -2093 1215
rect -2293 1165 -2277 1199
rect -2109 1165 -2093 1199
rect -2293 1118 -2093 1165
rect -2035 1199 -1835 1215
rect -2035 1165 -2019 1199
rect -1851 1165 -1835 1199
rect -2035 1118 -1835 1165
rect -1777 1199 -1577 1215
rect -1777 1165 -1761 1199
rect -1593 1165 -1577 1199
rect -1777 1118 -1577 1165
rect -1519 1199 -1319 1215
rect -1519 1165 -1503 1199
rect -1335 1165 -1319 1199
rect -1519 1118 -1319 1165
rect -1261 1199 -1061 1215
rect -1261 1165 -1245 1199
rect -1077 1165 -1061 1199
rect -1261 1118 -1061 1165
rect -1003 1199 -803 1215
rect -1003 1165 -987 1199
rect -819 1165 -803 1199
rect -1003 1118 -803 1165
rect -745 1199 -545 1215
rect -745 1165 -729 1199
rect -561 1165 -545 1199
rect -745 1118 -545 1165
rect -487 1199 -287 1215
rect -487 1165 -471 1199
rect -303 1165 -287 1199
rect -487 1118 -287 1165
rect -229 1199 -29 1215
rect -229 1165 -213 1199
rect -45 1165 -29 1199
rect -229 1118 -29 1165
rect 29 1199 229 1215
rect 29 1165 45 1199
rect 213 1165 229 1199
rect 29 1118 229 1165
rect 287 1199 487 1215
rect 287 1165 303 1199
rect 471 1165 487 1199
rect 287 1118 487 1165
rect 545 1199 745 1215
rect 545 1165 561 1199
rect 729 1165 745 1199
rect 545 1118 745 1165
rect 803 1199 1003 1215
rect 803 1165 819 1199
rect 987 1165 1003 1199
rect 803 1118 1003 1165
rect 1061 1199 1261 1215
rect 1061 1165 1077 1199
rect 1245 1165 1261 1199
rect 1061 1118 1261 1165
rect 1319 1199 1519 1215
rect 1319 1165 1335 1199
rect 1503 1165 1519 1199
rect 1319 1118 1519 1165
rect 1577 1199 1777 1215
rect 1577 1165 1593 1199
rect 1761 1165 1777 1199
rect 1577 1118 1777 1165
rect 1835 1199 2035 1215
rect 1835 1165 1851 1199
rect 2019 1165 2035 1199
rect 1835 1118 2035 1165
rect 2093 1199 2293 1215
rect 2093 1165 2109 1199
rect 2277 1165 2293 1199
rect 2093 1118 2293 1165
rect 2351 1199 2551 1215
rect 2351 1165 2367 1199
rect 2535 1165 2551 1199
rect 2351 1118 2551 1165
rect 2609 1199 2809 1215
rect 2609 1165 2625 1199
rect 2793 1165 2809 1199
rect 2609 1118 2809 1165
rect 2867 1199 3067 1215
rect 2867 1165 2883 1199
rect 3051 1165 3067 1199
rect 2867 1118 3067 1165
rect 3125 1199 3325 1215
rect 3125 1165 3141 1199
rect 3309 1165 3325 1199
rect 3125 1118 3325 1165
rect 3383 1199 3583 1215
rect 3383 1165 3399 1199
rect 3567 1165 3583 1199
rect 3383 1118 3583 1165
rect -3583 71 -3383 118
rect -3583 37 -3567 71
rect -3399 37 -3383 71
rect -3583 21 -3383 37
rect -3325 71 -3125 118
rect -3325 37 -3309 71
rect -3141 37 -3125 71
rect -3325 21 -3125 37
rect -3067 71 -2867 118
rect -3067 37 -3051 71
rect -2883 37 -2867 71
rect -3067 21 -2867 37
rect -2809 71 -2609 118
rect -2809 37 -2793 71
rect -2625 37 -2609 71
rect -2809 21 -2609 37
rect -2551 71 -2351 118
rect -2551 37 -2535 71
rect -2367 37 -2351 71
rect -2551 21 -2351 37
rect -2293 71 -2093 118
rect -2293 37 -2277 71
rect -2109 37 -2093 71
rect -2293 21 -2093 37
rect -2035 71 -1835 118
rect -2035 37 -2019 71
rect -1851 37 -1835 71
rect -2035 21 -1835 37
rect -1777 71 -1577 118
rect -1777 37 -1761 71
rect -1593 37 -1577 71
rect -1777 21 -1577 37
rect -1519 71 -1319 118
rect -1519 37 -1503 71
rect -1335 37 -1319 71
rect -1519 21 -1319 37
rect -1261 71 -1061 118
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1261 21 -1061 37
rect -1003 71 -803 118
rect -1003 37 -987 71
rect -819 37 -803 71
rect -1003 21 -803 37
rect -745 71 -545 118
rect -745 37 -729 71
rect -561 37 -545 71
rect -745 21 -545 37
rect -487 71 -287 118
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 118
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 118
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 118
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect 545 71 745 118
rect 545 37 561 71
rect 729 37 745 71
rect 545 21 745 37
rect 803 71 1003 118
rect 803 37 819 71
rect 987 37 1003 71
rect 803 21 1003 37
rect 1061 71 1261 118
rect 1061 37 1077 71
rect 1245 37 1261 71
rect 1061 21 1261 37
rect 1319 71 1519 118
rect 1319 37 1335 71
rect 1503 37 1519 71
rect 1319 21 1519 37
rect 1577 71 1777 118
rect 1577 37 1593 71
rect 1761 37 1777 71
rect 1577 21 1777 37
rect 1835 71 2035 118
rect 1835 37 1851 71
rect 2019 37 2035 71
rect 1835 21 2035 37
rect 2093 71 2293 118
rect 2093 37 2109 71
rect 2277 37 2293 71
rect 2093 21 2293 37
rect 2351 71 2551 118
rect 2351 37 2367 71
rect 2535 37 2551 71
rect 2351 21 2551 37
rect 2609 71 2809 118
rect 2609 37 2625 71
rect 2793 37 2809 71
rect 2609 21 2809 37
rect 2867 71 3067 118
rect 2867 37 2883 71
rect 3051 37 3067 71
rect 2867 21 3067 37
rect 3125 71 3325 118
rect 3125 37 3141 71
rect 3309 37 3325 71
rect 3125 21 3325 37
rect 3383 71 3583 118
rect 3383 37 3399 71
rect 3567 37 3583 71
rect 3383 21 3583 37
rect -3583 -37 -3383 -21
rect -3583 -71 -3567 -37
rect -3399 -71 -3383 -37
rect -3583 -118 -3383 -71
rect -3325 -37 -3125 -21
rect -3325 -71 -3309 -37
rect -3141 -71 -3125 -37
rect -3325 -118 -3125 -71
rect -3067 -37 -2867 -21
rect -3067 -71 -3051 -37
rect -2883 -71 -2867 -37
rect -3067 -118 -2867 -71
rect -2809 -37 -2609 -21
rect -2809 -71 -2793 -37
rect -2625 -71 -2609 -37
rect -2809 -118 -2609 -71
rect -2551 -37 -2351 -21
rect -2551 -71 -2535 -37
rect -2367 -71 -2351 -37
rect -2551 -118 -2351 -71
rect -2293 -37 -2093 -21
rect -2293 -71 -2277 -37
rect -2109 -71 -2093 -37
rect -2293 -118 -2093 -71
rect -2035 -37 -1835 -21
rect -2035 -71 -2019 -37
rect -1851 -71 -1835 -37
rect -2035 -118 -1835 -71
rect -1777 -37 -1577 -21
rect -1777 -71 -1761 -37
rect -1593 -71 -1577 -37
rect -1777 -118 -1577 -71
rect -1519 -37 -1319 -21
rect -1519 -71 -1503 -37
rect -1335 -71 -1319 -37
rect -1519 -118 -1319 -71
rect -1261 -37 -1061 -21
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1261 -118 -1061 -71
rect -1003 -37 -803 -21
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -1003 -118 -803 -71
rect -745 -37 -545 -21
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -745 -118 -545 -71
rect -487 -37 -287 -21
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -487 -118 -287 -71
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -118 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -118 229 -71
rect 287 -37 487 -21
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 287 -118 487 -71
rect 545 -37 745 -21
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 545 -118 745 -71
rect 803 -37 1003 -21
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 803 -118 1003 -71
rect 1061 -37 1261 -21
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect 1061 -118 1261 -71
rect 1319 -37 1519 -21
rect 1319 -71 1335 -37
rect 1503 -71 1519 -37
rect 1319 -118 1519 -71
rect 1577 -37 1777 -21
rect 1577 -71 1593 -37
rect 1761 -71 1777 -37
rect 1577 -118 1777 -71
rect 1835 -37 2035 -21
rect 1835 -71 1851 -37
rect 2019 -71 2035 -37
rect 1835 -118 2035 -71
rect 2093 -37 2293 -21
rect 2093 -71 2109 -37
rect 2277 -71 2293 -37
rect 2093 -118 2293 -71
rect 2351 -37 2551 -21
rect 2351 -71 2367 -37
rect 2535 -71 2551 -37
rect 2351 -118 2551 -71
rect 2609 -37 2809 -21
rect 2609 -71 2625 -37
rect 2793 -71 2809 -37
rect 2609 -118 2809 -71
rect 2867 -37 3067 -21
rect 2867 -71 2883 -37
rect 3051 -71 3067 -37
rect 2867 -118 3067 -71
rect 3125 -37 3325 -21
rect 3125 -71 3141 -37
rect 3309 -71 3325 -37
rect 3125 -118 3325 -71
rect 3383 -37 3583 -21
rect 3383 -71 3399 -37
rect 3567 -71 3583 -37
rect 3383 -118 3583 -71
rect -3583 -1165 -3383 -1118
rect -3583 -1199 -3567 -1165
rect -3399 -1199 -3383 -1165
rect -3583 -1215 -3383 -1199
rect -3325 -1165 -3125 -1118
rect -3325 -1199 -3309 -1165
rect -3141 -1199 -3125 -1165
rect -3325 -1215 -3125 -1199
rect -3067 -1165 -2867 -1118
rect -3067 -1199 -3051 -1165
rect -2883 -1199 -2867 -1165
rect -3067 -1215 -2867 -1199
rect -2809 -1165 -2609 -1118
rect -2809 -1199 -2793 -1165
rect -2625 -1199 -2609 -1165
rect -2809 -1215 -2609 -1199
rect -2551 -1165 -2351 -1118
rect -2551 -1199 -2535 -1165
rect -2367 -1199 -2351 -1165
rect -2551 -1215 -2351 -1199
rect -2293 -1165 -2093 -1118
rect -2293 -1199 -2277 -1165
rect -2109 -1199 -2093 -1165
rect -2293 -1215 -2093 -1199
rect -2035 -1165 -1835 -1118
rect -2035 -1199 -2019 -1165
rect -1851 -1199 -1835 -1165
rect -2035 -1215 -1835 -1199
rect -1777 -1165 -1577 -1118
rect -1777 -1199 -1761 -1165
rect -1593 -1199 -1577 -1165
rect -1777 -1215 -1577 -1199
rect -1519 -1165 -1319 -1118
rect -1519 -1199 -1503 -1165
rect -1335 -1199 -1319 -1165
rect -1519 -1215 -1319 -1199
rect -1261 -1165 -1061 -1118
rect -1261 -1199 -1245 -1165
rect -1077 -1199 -1061 -1165
rect -1261 -1215 -1061 -1199
rect -1003 -1165 -803 -1118
rect -1003 -1199 -987 -1165
rect -819 -1199 -803 -1165
rect -1003 -1215 -803 -1199
rect -745 -1165 -545 -1118
rect -745 -1199 -729 -1165
rect -561 -1199 -545 -1165
rect -745 -1215 -545 -1199
rect -487 -1165 -287 -1118
rect -487 -1199 -471 -1165
rect -303 -1199 -287 -1165
rect -487 -1215 -287 -1199
rect -229 -1165 -29 -1118
rect -229 -1199 -213 -1165
rect -45 -1199 -29 -1165
rect -229 -1215 -29 -1199
rect 29 -1165 229 -1118
rect 29 -1199 45 -1165
rect 213 -1199 229 -1165
rect 29 -1215 229 -1199
rect 287 -1165 487 -1118
rect 287 -1199 303 -1165
rect 471 -1199 487 -1165
rect 287 -1215 487 -1199
rect 545 -1165 745 -1118
rect 545 -1199 561 -1165
rect 729 -1199 745 -1165
rect 545 -1215 745 -1199
rect 803 -1165 1003 -1118
rect 803 -1199 819 -1165
rect 987 -1199 1003 -1165
rect 803 -1215 1003 -1199
rect 1061 -1165 1261 -1118
rect 1061 -1199 1077 -1165
rect 1245 -1199 1261 -1165
rect 1061 -1215 1261 -1199
rect 1319 -1165 1519 -1118
rect 1319 -1199 1335 -1165
rect 1503 -1199 1519 -1165
rect 1319 -1215 1519 -1199
rect 1577 -1165 1777 -1118
rect 1577 -1199 1593 -1165
rect 1761 -1199 1777 -1165
rect 1577 -1215 1777 -1199
rect 1835 -1165 2035 -1118
rect 1835 -1199 1851 -1165
rect 2019 -1199 2035 -1165
rect 1835 -1215 2035 -1199
rect 2093 -1165 2293 -1118
rect 2093 -1199 2109 -1165
rect 2277 -1199 2293 -1165
rect 2093 -1215 2293 -1199
rect 2351 -1165 2551 -1118
rect 2351 -1199 2367 -1165
rect 2535 -1199 2551 -1165
rect 2351 -1215 2551 -1199
rect 2609 -1165 2809 -1118
rect 2609 -1199 2625 -1165
rect 2793 -1199 2809 -1165
rect 2609 -1215 2809 -1199
rect 2867 -1165 3067 -1118
rect 2867 -1199 2883 -1165
rect 3051 -1199 3067 -1165
rect 2867 -1215 3067 -1199
rect 3125 -1165 3325 -1118
rect 3125 -1199 3141 -1165
rect 3309 -1199 3325 -1165
rect 3125 -1215 3325 -1199
rect 3383 -1165 3583 -1118
rect 3383 -1199 3399 -1165
rect 3567 -1199 3583 -1165
rect 3383 -1215 3583 -1199
rect -3583 -1273 -3383 -1257
rect -3583 -1307 -3567 -1273
rect -3399 -1307 -3383 -1273
rect -3583 -1354 -3383 -1307
rect -3325 -1273 -3125 -1257
rect -3325 -1307 -3309 -1273
rect -3141 -1307 -3125 -1273
rect -3325 -1354 -3125 -1307
rect -3067 -1273 -2867 -1257
rect -3067 -1307 -3051 -1273
rect -2883 -1307 -2867 -1273
rect -3067 -1354 -2867 -1307
rect -2809 -1273 -2609 -1257
rect -2809 -1307 -2793 -1273
rect -2625 -1307 -2609 -1273
rect -2809 -1354 -2609 -1307
rect -2551 -1273 -2351 -1257
rect -2551 -1307 -2535 -1273
rect -2367 -1307 -2351 -1273
rect -2551 -1354 -2351 -1307
rect -2293 -1273 -2093 -1257
rect -2293 -1307 -2277 -1273
rect -2109 -1307 -2093 -1273
rect -2293 -1354 -2093 -1307
rect -2035 -1273 -1835 -1257
rect -2035 -1307 -2019 -1273
rect -1851 -1307 -1835 -1273
rect -2035 -1354 -1835 -1307
rect -1777 -1273 -1577 -1257
rect -1777 -1307 -1761 -1273
rect -1593 -1307 -1577 -1273
rect -1777 -1354 -1577 -1307
rect -1519 -1273 -1319 -1257
rect -1519 -1307 -1503 -1273
rect -1335 -1307 -1319 -1273
rect -1519 -1354 -1319 -1307
rect -1261 -1273 -1061 -1257
rect -1261 -1307 -1245 -1273
rect -1077 -1307 -1061 -1273
rect -1261 -1354 -1061 -1307
rect -1003 -1273 -803 -1257
rect -1003 -1307 -987 -1273
rect -819 -1307 -803 -1273
rect -1003 -1354 -803 -1307
rect -745 -1273 -545 -1257
rect -745 -1307 -729 -1273
rect -561 -1307 -545 -1273
rect -745 -1354 -545 -1307
rect -487 -1273 -287 -1257
rect -487 -1307 -471 -1273
rect -303 -1307 -287 -1273
rect -487 -1354 -287 -1307
rect -229 -1273 -29 -1257
rect -229 -1307 -213 -1273
rect -45 -1307 -29 -1273
rect -229 -1354 -29 -1307
rect 29 -1273 229 -1257
rect 29 -1307 45 -1273
rect 213 -1307 229 -1273
rect 29 -1354 229 -1307
rect 287 -1273 487 -1257
rect 287 -1307 303 -1273
rect 471 -1307 487 -1273
rect 287 -1354 487 -1307
rect 545 -1273 745 -1257
rect 545 -1307 561 -1273
rect 729 -1307 745 -1273
rect 545 -1354 745 -1307
rect 803 -1273 1003 -1257
rect 803 -1307 819 -1273
rect 987 -1307 1003 -1273
rect 803 -1354 1003 -1307
rect 1061 -1273 1261 -1257
rect 1061 -1307 1077 -1273
rect 1245 -1307 1261 -1273
rect 1061 -1354 1261 -1307
rect 1319 -1273 1519 -1257
rect 1319 -1307 1335 -1273
rect 1503 -1307 1519 -1273
rect 1319 -1354 1519 -1307
rect 1577 -1273 1777 -1257
rect 1577 -1307 1593 -1273
rect 1761 -1307 1777 -1273
rect 1577 -1354 1777 -1307
rect 1835 -1273 2035 -1257
rect 1835 -1307 1851 -1273
rect 2019 -1307 2035 -1273
rect 1835 -1354 2035 -1307
rect 2093 -1273 2293 -1257
rect 2093 -1307 2109 -1273
rect 2277 -1307 2293 -1273
rect 2093 -1354 2293 -1307
rect 2351 -1273 2551 -1257
rect 2351 -1307 2367 -1273
rect 2535 -1307 2551 -1273
rect 2351 -1354 2551 -1307
rect 2609 -1273 2809 -1257
rect 2609 -1307 2625 -1273
rect 2793 -1307 2809 -1273
rect 2609 -1354 2809 -1307
rect 2867 -1273 3067 -1257
rect 2867 -1307 2883 -1273
rect 3051 -1307 3067 -1273
rect 2867 -1354 3067 -1307
rect 3125 -1273 3325 -1257
rect 3125 -1307 3141 -1273
rect 3309 -1307 3325 -1273
rect 3125 -1354 3325 -1307
rect 3383 -1273 3583 -1257
rect 3383 -1307 3399 -1273
rect 3567 -1307 3583 -1273
rect 3383 -1354 3583 -1307
rect -3583 -2401 -3383 -2354
rect -3583 -2435 -3567 -2401
rect -3399 -2435 -3383 -2401
rect -3583 -2451 -3383 -2435
rect -3325 -2401 -3125 -2354
rect -3325 -2435 -3309 -2401
rect -3141 -2435 -3125 -2401
rect -3325 -2451 -3125 -2435
rect -3067 -2401 -2867 -2354
rect -3067 -2435 -3051 -2401
rect -2883 -2435 -2867 -2401
rect -3067 -2451 -2867 -2435
rect -2809 -2401 -2609 -2354
rect -2809 -2435 -2793 -2401
rect -2625 -2435 -2609 -2401
rect -2809 -2451 -2609 -2435
rect -2551 -2401 -2351 -2354
rect -2551 -2435 -2535 -2401
rect -2367 -2435 -2351 -2401
rect -2551 -2451 -2351 -2435
rect -2293 -2401 -2093 -2354
rect -2293 -2435 -2277 -2401
rect -2109 -2435 -2093 -2401
rect -2293 -2451 -2093 -2435
rect -2035 -2401 -1835 -2354
rect -2035 -2435 -2019 -2401
rect -1851 -2435 -1835 -2401
rect -2035 -2451 -1835 -2435
rect -1777 -2401 -1577 -2354
rect -1777 -2435 -1761 -2401
rect -1593 -2435 -1577 -2401
rect -1777 -2451 -1577 -2435
rect -1519 -2401 -1319 -2354
rect -1519 -2435 -1503 -2401
rect -1335 -2435 -1319 -2401
rect -1519 -2451 -1319 -2435
rect -1261 -2401 -1061 -2354
rect -1261 -2435 -1245 -2401
rect -1077 -2435 -1061 -2401
rect -1261 -2451 -1061 -2435
rect -1003 -2401 -803 -2354
rect -1003 -2435 -987 -2401
rect -819 -2435 -803 -2401
rect -1003 -2451 -803 -2435
rect -745 -2401 -545 -2354
rect -745 -2435 -729 -2401
rect -561 -2435 -545 -2401
rect -745 -2451 -545 -2435
rect -487 -2401 -287 -2354
rect -487 -2435 -471 -2401
rect -303 -2435 -287 -2401
rect -487 -2451 -287 -2435
rect -229 -2401 -29 -2354
rect -229 -2435 -213 -2401
rect -45 -2435 -29 -2401
rect -229 -2451 -29 -2435
rect 29 -2401 229 -2354
rect 29 -2435 45 -2401
rect 213 -2435 229 -2401
rect 29 -2451 229 -2435
rect 287 -2401 487 -2354
rect 287 -2435 303 -2401
rect 471 -2435 487 -2401
rect 287 -2451 487 -2435
rect 545 -2401 745 -2354
rect 545 -2435 561 -2401
rect 729 -2435 745 -2401
rect 545 -2451 745 -2435
rect 803 -2401 1003 -2354
rect 803 -2435 819 -2401
rect 987 -2435 1003 -2401
rect 803 -2451 1003 -2435
rect 1061 -2401 1261 -2354
rect 1061 -2435 1077 -2401
rect 1245 -2435 1261 -2401
rect 1061 -2451 1261 -2435
rect 1319 -2401 1519 -2354
rect 1319 -2435 1335 -2401
rect 1503 -2435 1519 -2401
rect 1319 -2451 1519 -2435
rect 1577 -2401 1777 -2354
rect 1577 -2435 1593 -2401
rect 1761 -2435 1777 -2401
rect 1577 -2451 1777 -2435
rect 1835 -2401 2035 -2354
rect 1835 -2435 1851 -2401
rect 2019 -2435 2035 -2401
rect 1835 -2451 2035 -2435
rect 2093 -2401 2293 -2354
rect 2093 -2435 2109 -2401
rect 2277 -2435 2293 -2401
rect 2093 -2451 2293 -2435
rect 2351 -2401 2551 -2354
rect 2351 -2435 2367 -2401
rect 2535 -2435 2551 -2401
rect 2351 -2451 2551 -2435
rect 2609 -2401 2809 -2354
rect 2609 -2435 2625 -2401
rect 2793 -2435 2809 -2401
rect 2609 -2451 2809 -2435
rect 2867 -2401 3067 -2354
rect 2867 -2435 2883 -2401
rect 3051 -2435 3067 -2401
rect 2867 -2451 3067 -2435
rect 3125 -2401 3325 -2354
rect 3125 -2435 3141 -2401
rect 3309 -2435 3325 -2401
rect 3125 -2451 3325 -2435
rect 3383 -2401 3583 -2354
rect 3383 -2435 3399 -2401
rect 3567 -2435 3583 -2401
rect 3383 -2451 3583 -2435
<< polycont >>
rect -3567 2401 -3399 2435
rect -3309 2401 -3141 2435
rect -3051 2401 -2883 2435
rect -2793 2401 -2625 2435
rect -2535 2401 -2367 2435
rect -2277 2401 -2109 2435
rect -2019 2401 -1851 2435
rect -1761 2401 -1593 2435
rect -1503 2401 -1335 2435
rect -1245 2401 -1077 2435
rect -987 2401 -819 2435
rect -729 2401 -561 2435
rect -471 2401 -303 2435
rect -213 2401 -45 2435
rect 45 2401 213 2435
rect 303 2401 471 2435
rect 561 2401 729 2435
rect 819 2401 987 2435
rect 1077 2401 1245 2435
rect 1335 2401 1503 2435
rect 1593 2401 1761 2435
rect 1851 2401 2019 2435
rect 2109 2401 2277 2435
rect 2367 2401 2535 2435
rect 2625 2401 2793 2435
rect 2883 2401 3051 2435
rect 3141 2401 3309 2435
rect 3399 2401 3567 2435
rect -3567 1273 -3399 1307
rect -3309 1273 -3141 1307
rect -3051 1273 -2883 1307
rect -2793 1273 -2625 1307
rect -2535 1273 -2367 1307
rect -2277 1273 -2109 1307
rect -2019 1273 -1851 1307
rect -1761 1273 -1593 1307
rect -1503 1273 -1335 1307
rect -1245 1273 -1077 1307
rect -987 1273 -819 1307
rect -729 1273 -561 1307
rect -471 1273 -303 1307
rect -213 1273 -45 1307
rect 45 1273 213 1307
rect 303 1273 471 1307
rect 561 1273 729 1307
rect 819 1273 987 1307
rect 1077 1273 1245 1307
rect 1335 1273 1503 1307
rect 1593 1273 1761 1307
rect 1851 1273 2019 1307
rect 2109 1273 2277 1307
rect 2367 1273 2535 1307
rect 2625 1273 2793 1307
rect 2883 1273 3051 1307
rect 3141 1273 3309 1307
rect 3399 1273 3567 1307
rect -3567 1165 -3399 1199
rect -3309 1165 -3141 1199
rect -3051 1165 -2883 1199
rect -2793 1165 -2625 1199
rect -2535 1165 -2367 1199
rect -2277 1165 -2109 1199
rect -2019 1165 -1851 1199
rect -1761 1165 -1593 1199
rect -1503 1165 -1335 1199
rect -1245 1165 -1077 1199
rect -987 1165 -819 1199
rect -729 1165 -561 1199
rect -471 1165 -303 1199
rect -213 1165 -45 1199
rect 45 1165 213 1199
rect 303 1165 471 1199
rect 561 1165 729 1199
rect 819 1165 987 1199
rect 1077 1165 1245 1199
rect 1335 1165 1503 1199
rect 1593 1165 1761 1199
rect 1851 1165 2019 1199
rect 2109 1165 2277 1199
rect 2367 1165 2535 1199
rect 2625 1165 2793 1199
rect 2883 1165 3051 1199
rect 3141 1165 3309 1199
rect 3399 1165 3567 1199
rect -3567 37 -3399 71
rect -3309 37 -3141 71
rect -3051 37 -2883 71
rect -2793 37 -2625 71
rect -2535 37 -2367 71
rect -2277 37 -2109 71
rect -2019 37 -1851 71
rect -1761 37 -1593 71
rect -1503 37 -1335 71
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect 1335 37 1503 71
rect 1593 37 1761 71
rect 1851 37 2019 71
rect 2109 37 2277 71
rect 2367 37 2535 71
rect 2625 37 2793 71
rect 2883 37 3051 71
rect 3141 37 3309 71
rect 3399 37 3567 71
rect -3567 -71 -3399 -37
rect -3309 -71 -3141 -37
rect -3051 -71 -2883 -37
rect -2793 -71 -2625 -37
rect -2535 -71 -2367 -37
rect -2277 -71 -2109 -37
rect -2019 -71 -1851 -37
rect -1761 -71 -1593 -37
rect -1503 -71 -1335 -37
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect 1335 -71 1503 -37
rect 1593 -71 1761 -37
rect 1851 -71 2019 -37
rect 2109 -71 2277 -37
rect 2367 -71 2535 -37
rect 2625 -71 2793 -37
rect 2883 -71 3051 -37
rect 3141 -71 3309 -37
rect 3399 -71 3567 -37
rect -3567 -1199 -3399 -1165
rect -3309 -1199 -3141 -1165
rect -3051 -1199 -2883 -1165
rect -2793 -1199 -2625 -1165
rect -2535 -1199 -2367 -1165
rect -2277 -1199 -2109 -1165
rect -2019 -1199 -1851 -1165
rect -1761 -1199 -1593 -1165
rect -1503 -1199 -1335 -1165
rect -1245 -1199 -1077 -1165
rect -987 -1199 -819 -1165
rect -729 -1199 -561 -1165
rect -471 -1199 -303 -1165
rect -213 -1199 -45 -1165
rect 45 -1199 213 -1165
rect 303 -1199 471 -1165
rect 561 -1199 729 -1165
rect 819 -1199 987 -1165
rect 1077 -1199 1245 -1165
rect 1335 -1199 1503 -1165
rect 1593 -1199 1761 -1165
rect 1851 -1199 2019 -1165
rect 2109 -1199 2277 -1165
rect 2367 -1199 2535 -1165
rect 2625 -1199 2793 -1165
rect 2883 -1199 3051 -1165
rect 3141 -1199 3309 -1165
rect 3399 -1199 3567 -1165
rect -3567 -1307 -3399 -1273
rect -3309 -1307 -3141 -1273
rect -3051 -1307 -2883 -1273
rect -2793 -1307 -2625 -1273
rect -2535 -1307 -2367 -1273
rect -2277 -1307 -2109 -1273
rect -2019 -1307 -1851 -1273
rect -1761 -1307 -1593 -1273
rect -1503 -1307 -1335 -1273
rect -1245 -1307 -1077 -1273
rect -987 -1307 -819 -1273
rect -729 -1307 -561 -1273
rect -471 -1307 -303 -1273
rect -213 -1307 -45 -1273
rect 45 -1307 213 -1273
rect 303 -1307 471 -1273
rect 561 -1307 729 -1273
rect 819 -1307 987 -1273
rect 1077 -1307 1245 -1273
rect 1335 -1307 1503 -1273
rect 1593 -1307 1761 -1273
rect 1851 -1307 2019 -1273
rect 2109 -1307 2277 -1273
rect 2367 -1307 2535 -1273
rect 2625 -1307 2793 -1273
rect 2883 -1307 3051 -1273
rect 3141 -1307 3309 -1273
rect 3399 -1307 3567 -1273
rect -3567 -2435 -3399 -2401
rect -3309 -2435 -3141 -2401
rect -3051 -2435 -2883 -2401
rect -2793 -2435 -2625 -2401
rect -2535 -2435 -2367 -2401
rect -2277 -2435 -2109 -2401
rect -2019 -2435 -1851 -2401
rect -1761 -2435 -1593 -2401
rect -1503 -2435 -1335 -2401
rect -1245 -2435 -1077 -2401
rect -987 -2435 -819 -2401
rect -729 -2435 -561 -2401
rect -471 -2435 -303 -2401
rect -213 -2435 -45 -2401
rect 45 -2435 213 -2401
rect 303 -2435 471 -2401
rect 561 -2435 729 -2401
rect 819 -2435 987 -2401
rect 1077 -2435 1245 -2401
rect 1335 -2435 1503 -2401
rect 1593 -2435 1761 -2401
rect 1851 -2435 2019 -2401
rect 2109 -2435 2277 -2401
rect 2367 -2435 2535 -2401
rect 2625 -2435 2793 -2401
rect 2883 -2435 3051 -2401
rect 3141 -2435 3309 -2401
rect 3399 -2435 3567 -2401
<< locali >>
rect -3763 2539 -3667 2573
rect 3667 2539 3763 2573
rect -3763 2477 -3729 2539
rect 3729 2477 3763 2539
rect -3583 2401 -3567 2435
rect -3399 2401 -3383 2435
rect -3325 2401 -3309 2435
rect -3141 2401 -3125 2435
rect -3067 2401 -3051 2435
rect -2883 2401 -2867 2435
rect -2809 2401 -2793 2435
rect -2625 2401 -2609 2435
rect -2551 2401 -2535 2435
rect -2367 2401 -2351 2435
rect -2293 2401 -2277 2435
rect -2109 2401 -2093 2435
rect -2035 2401 -2019 2435
rect -1851 2401 -1835 2435
rect -1777 2401 -1761 2435
rect -1593 2401 -1577 2435
rect -1519 2401 -1503 2435
rect -1335 2401 -1319 2435
rect -1261 2401 -1245 2435
rect -1077 2401 -1061 2435
rect -1003 2401 -987 2435
rect -819 2401 -803 2435
rect -745 2401 -729 2435
rect -561 2401 -545 2435
rect -487 2401 -471 2435
rect -303 2401 -287 2435
rect -229 2401 -213 2435
rect -45 2401 -29 2435
rect 29 2401 45 2435
rect 213 2401 229 2435
rect 287 2401 303 2435
rect 471 2401 487 2435
rect 545 2401 561 2435
rect 729 2401 745 2435
rect 803 2401 819 2435
rect 987 2401 1003 2435
rect 1061 2401 1077 2435
rect 1245 2401 1261 2435
rect 1319 2401 1335 2435
rect 1503 2401 1519 2435
rect 1577 2401 1593 2435
rect 1761 2401 1777 2435
rect 1835 2401 1851 2435
rect 2019 2401 2035 2435
rect 2093 2401 2109 2435
rect 2277 2401 2293 2435
rect 2351 2401 2367 2435
rect 2535 2401 2551 2435
rect 2609 2401 2625 2435
rect 2793 2401 2809 2435
rect 2867 2401 2883 2435
rect 3051 2401 3067 2435
rect 3125 2401 3141 2435
rect 3309 2401 3325 2435
rect 3383 2401 3399 2435
rect 3567 2401 3583 2435
rect -3629 2342 -3595 2358
rect -3629 1350 -3595 1366
rect -3371 2342 -3337 2358
rect -3371 1350 -3337 1366
rect -3113 2342 -3079 2358
rect -3113 1350 -3079 1366
rect -2855 2342 -2821 2358
rect -2855 1350 -2821 1366
rect -2597 2342 -2563 2358
rect -2597 1350 -2563 1366
rect -2339 2342 -2305 2358
rect -2339 1350 -2305 1366
rect -2081 2342 -2047 2358
rect -2081 1350 -2047 1366
rect -1823 2342 -1789 2358
rect -1823 1350 -1789 1366
rect -1565 2342 -1531 2358
rect -1565 1350 -1531 1366
rect -1307 2342 -1273 2358
rect -1307 1350 -1273 1366
rect -1049 2342 -1015 2358
rect -1049 1350 -1015 1366
rect -791 2342 -757 2358
rect -791 1350 -757 1366
rect -533 2342 -499 2358
rect -533 1350 -499 1366
rect -275 2342 -241 2358
rect -275 1350 -241 1366
rect -17 2342 17 2358
rect -17 1350 17 1366
rect 241 2342 275 2358
rect 241 1350 275 1366
rect 499 2342 533 2358
rect 499 1350 533 1366
rect 757 2342 791 2358
rect 757 1350 791 1366
rect 1015 2342 1049 2358
rect 1015 1350 1049 1366
rect 1273 2342 1307 2358
rect 1273 1350 1307 1366
rect 1531 2342 1565 2358
rect 1531 1350 1565 1366
rect 1789 2342 1823 2358
rect 1789 1350 1823 1366
rect 2047 2342 2081 2358
rect 2047 1350 2081 1366
rect 2305 2342 2339 2358
rect 2305 1350 2339 1366
rect 2563 2342 2597 2358
rect 2563 1350 2597 1366
rect 2821 2342 2855 2358
rect 2821 1350 2855 1366
rect 3079 2342 3113 2358
rect 3079 1350 3113 1366
rect 3337 2342 3371 2358
rect 3337 1350 3371 1366
rect 3595 2342 3629 2358
rect 3595 1350 3629 1366
rect -3583 1273 -3567 1307
rect -3399 1273 -3383 1307
rect -3325 1273 -3309 1307
rect -3141 1273 -3125 1307
rect -3067 1273 -3051 1307
rect -2883 1273 -2867 1307
rect -2809 1273 -2793 1307
rect -2625 1273 -2609 1307
rect -2551 1273 -2535 1307
rect -2367 1273 -2351 1307
rect -2293 1273 -2277 1307
rect -2109 1273 -2093 1307
rect -2035 1273 -2019 1307
rect -1851 1273 -1835 1307
rect -1777 1273 -1761 1307
rect -1593 1273 -1577 1307
rect -1519 1273 -1503 1307
rect -1335 1273 -1319 1307
rect -1261 1273 -1245 1307
rect -1077 1273 -1061 1307
rect -1003 1273 -987 1307
rect -819 1273 -803 1307
rect -745 1273 -729 1307
rect -561 1273 -545 1307
rect -487 1273 -471 1307
rect -303 1273 -287 1307
rect -229 1273 -213 1307
rect -45 1273 -29 1307
rect 29 1273 45 1307
rect 213 1273 229 1307
rect 287 1273 303 1307
rect 471 1273 487 1307
rect 545 1273 561 1307
rect 729 1273 745 1307
rect 803 1273 819 1307
rect 987 1273 1003 1307
rect 1061 1273 1077 1307
rect 1245 1273 1261 1307
rect 1319 1273 1335 1307
rect 1503 1273 1519 1307
rect 1577 1273 1593 1307
rect 1761 1273 1777 1307
rect 1835 1273 1851 1307
rect 2019 1273 2035 1307
rect 2093 1273 2109 1307
rect 2277 1273 2293 1307
rect 2351 1273 2367 1307
rect 2535 1273 2551 1307
rect 2609 1273 2625 1307
rect 2793 1273 2809 1307
rect 2867 1273 2883 1307
rect 3051 1273 3067 1307
rect 3125 1273 3141 1307
rect 3309 1273 3325 1307
rect 3383 1273 3399 1307
rect 3567 1273 3583 1307
rect -3583 1165 -3567 1199
rect -3399 1165 -3383 1199
rect -3325 1165 -3309 1199
rect -3141 1165 -3125 1199
rect -3067 1165 -3051 1199
rect -2883 1165 -2867 1199
rect -2809 1165 -2793 1199
rect -2625 1165 -2609 1199
rect -2551 1165 -2535 1199
rect -2367 1165 -2351 1199
rect -2293 1165 -2277 1199
rect -2109 1165 -2093 1199
rect -2035 1165 -2019 1199
rect -1851 1165 -1835 1199
rect -1777 1165 -1761 1199
rect -1593 1165 -1577 1199
rect -1519 1165 -1503 1199
rect -1335 1165 -1319 1199
rect -1261 1165 -1245 1199
rect -1077 1165 -1061 1199
rect -1003 1165 -987 1199
rect -819 1165 -803 1199
rect -745 1165 -729 1199
rect -561 1165 -545 1199
rect -487 1165 -471 1199
rect -303 1165 -287 1199
rect -229 1165 -213 1199
rect -45 1165 -29 1199
rect 29 1165 45 1199
rect 213 1165 229 1199
rect 287 1165 303 1199
rect 471 1165 487 1199
rect 545 1165 561 1199
rect 729 1165 745 1199
rect 803 1165 819 1199
rect 987 1165 1003 1199
rect 1061 1165 1077 1199
rect 1245 1165 1261 1199
rect 1319 1165 1335 1199
rect 1503 1165 1519 1199
rect 1577 1165 1593 1199
rect 1761 1165 1777 1199
rect 1835 1165 1851 1199
rect 2019 1165 2035 1199
rect 2093 1165 2109 1199
rect 2277 1165 2293 1199
rect 2351 1165 2367 1199
rect 2535 1165 2551 1199
rect 2609 1165 2625 1199
rect 2793 1165 2809 1199
rect 2867 1165 2883 1199
rect 3051 1165 3067 1199
rect 3125 1165 3141 1199
rect 3309 1165 3325 1199
rect 3383 1165 3399 1199
rect 3567 1165 3583 1199
rect -3629 1106 -3595 1122
rect -3629 114 -3595 130
rect -3371 1106 -3337 1122
rect -3371 114 -3337 130
rect -3113 1106 -3079 1122
rect -3113 114 -3079 130
rect -2855 1106 -2821 1122
rect -2855 114 -2821 130
rect -2597 1106 -2563 1122
rect -2597 114 -2563 130
rect -2339 1106 -2305 1122
rect -2339 114 -2305 130
rect -2081 1106 -2047 1122
rect -2081 114 -2047 130
rect -1823 1106 -1789 1122
rect -1823 114 -1789 130
rect -1565 1106 -1531 1122
rect -1565 114 -1531 130
rect -1307 1106 -1273 1122
rect -1307 114 -1273 130
rect -1049 1106 -1015 1122
rect -1049 114 -1015 130
rect -791 1106 -757 1122
rect -791 114 -757 130
rect -533 1106 -499 1122
rect -533 114 -499 130
rect -275 1106 -241 1122
rect -275 114 -241 130
rect -17 1106 17 1122
rect -17 114 17 130
rect 241 1106 275 1122
rect 241 114 275 130
rect 499 1106 533 1122
rect 499 114 533 130
rect 757 1106 791 1122
rect 757 114 791 130
rect 1015 1106 1049 1122
rect 1015 114 1049 130
rect 1273 1106 1307 1122
rect 1273 114 1307 130
rect 1531 1106 1565 1122
rect 1531 114 1565 130
rect 1789 1106 1823 1122
rect 1789 114 1823 130
rect 2047 1106 2081 1122
rect 2047 114 2081 130
rect 2305 1106 2339 1122
rect 2305 114 2339 130
rect 2563 1106 2597 1122
rect 2563 114 2597 130
rect 2821 1106 2855 1122
rect 2821 114 2855 130
rect 3079 1106 3113 1122
rect 3079 114 3113 130
rect 3337 1106 3371 1122
rect 3337 114 3371 130
rect 3595 1106 3629 1122
rect 3595 114 3629 130
rect -3583 37 -3567 71
rect -3399 37 -3383 71
rect -3325 37 -3309 71
rect -3141 37 -3125 71
rect -3067 37 -3051 71
rect -2883 37 -2867 71
rect -2809 37 -2793 71
rect -2625 37 -2609 71
rect -2551 37 -2535 71
rect -2367 37 -2351 71
rect -2293 37 -2277 71
rect -2109 37 -2093 71
rect -2035 37 -2019 71
rect -1851 37 -1835 71
rect -1777 37 -1761 71
rect -1593 37 -1577 71
rect -1519 37 -1503 71
rect -1335 37 -1319 71
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1003 37 -987 71
rect -819 37 -803 71
rect -745 37 -729 71
rect -561 37 -545 71
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect 545 37 561 71
rect 729 37 745 71
rect 803 37 819 71
rect 987 37 1003 71
rect 1061 37 1077 71
rect 1245 37 1261 71
rect 1319 37 1335 71
rect 1503 37 1519 71
rect 1577 37 1593 71
rect 1761 37 1777 71
rect 1835 37 1851 71
rect 2019 37 2035 71
rect 2093 37 2109 71
rect 2277 37 2293 71
rect 2351 37 2367 71
rect 2535 37 2551 71
rect 2609 37 2625 71
rect 2793 37 2809 71
rect 2867 37 2883 71
rect 3051 37 3067 71
rect 3125 37 3141 71
rect 3309 37 3325 71
rect 3383 37 3399 71
rect 3567 37 3583 71
rect -3583 -71 -3567 -37
rect -3399 -71 -3383 -37
rect -3325 -71 -3309 -37
rect -3141 -71 -3125 -37
rect -3067 -71 -3051 -37
rect -2883 -71 -2867 -37
rect -2809 -71 -2793 -37
rect -2625 -71 -2609 -37
rect -2551 -71 -2535 -37
rect -2367 -71 -2351 -37
rect -2293 -71 -2277 -37
rect -2109 -71 -2093 -37
rect -2035 -71 -2019 -37
rect -1851 -71 -1835 -37
rect -1777 -71 -1761 -37
rect -1593 -71 -1577 -37
rect -1519 -71 -1503 -37
rect -1335 -71 -1319 -37
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect 1319 -71 1335 -37
rect 1503 -71 1519 -37
rect 1577 -71 1593 -37
rect 1761 -71 1777 -37
rect 1835 -71 1851 -37
rect 2019 -71 2035 -37
rect 2093 -71 2109 -37
rect 2277 -71 2293 -37
rect 2351 -71 2367 -37
rect 2535 -71 2551 -37
rect 2609 -71 2625 -37
rect 2793 -71 2809 -37
rect 2867 -71 2883 -37
rect 3051 -71 3067 -37
rect 3125 -71 3141 -37
rect 3309 -71 3325 -37
rect 3383 -71 3399 -37
rect 3567 -71 3583 -37
rect -3629 -130 -3595 -114
rect -3629 -1122 -3595 -1106
rect -3371 -130 -3337 -114
rect -3371 -1122 -3337 -1106
rect -3113 -130 -3079 -114
rect -3113 -1122 -3079 -1106
rect -2855 -130 -2821 -114
rect -2855 -1122 -2821 -1106
rect -2597 -130 -2563 -114
rect -2597 -1122 -2563 -1106
rect -2339 -130 -2305 -114
rect -2339 -1122 -2305 -1106
rect -2081 -130 -2047 -114
rect -2081 -1122 -2047 -1106
rect -1823 -130 -1789 -114
rect -1823 -1122 -1789 -1106
rect -1565 -130 -1531 -114
rect -1565 -1122 -1531 -1106
rect -1307 -130 -1273 -114
rect -1307 -1122 -1273 -1106
rect -1049 -130 -1015 -114
rect -1049 -1122 -1015 -1106
rect -791 -130 -757 -114
rect -791 -1122 -757 -1106
rect -533 -130 -499 -114
rect -533 -1122 -499 -1106
rect -275 -130 -241 -114
rect -275 -1122 -241 -1106
rect -17 -130 17 -114
rect -17 -1122 17 -1106
rect 241 -130 275 -114
rect 241 -1122 275 -1106
rect 499 -130 533 -114
rect 499 -1122 533 -1106
rect 757 -130 791 -114
rect 757 -1122 791 -1106
rect 1015 -130 1049 -114
rect 1015 -1122 1049 -1106
rect 1273 -130 1307 -114
rect 1273 -1122 1307 -1106
rect 1531 -130 1565 -114
rect 1531 -1122 1565 -1106
rect 1789 -130 1823 -114
rect 1789 -1122 1823 -1106
rect 2047 -130 2081 -114
rect 2047 -1122 2081 -1106
rect 2305 -130 2339 -114
rect 2305 -1122 2339 -1106
rect 2563 -130 2597 -114
rect 2563 -1122 2597 -1106
rect 2821 -130 2855 -114
rect 2821 -1122 2855 -1106
rect 3079 -130 3113 -114
rect 3079 -1122 3113 -1106
rect 3337 -130 3371 -114
rect 3337 -1122 3371 -1106
rect 3595 -130 3629 -114
rect 3595 -1122 3629 -1106
rect -3583 -1199 -3567 -1165
rect -3399 -1199 -3383 -1165
rect -3325 -1199 -3309 -1165
rect -3141 -1199 -3125 -1165
rect -3067 -1199 -3051 -1165
rect -2883 -1199 -2867 -1165
rect -2809 -1199 -2793 -1165
rect -2625 -1199 -2609 -1165
rect -2551 -1199 -2535 -1165
rect -2367 -1199 -2351 -1165
rect -2293 -1199 -2277 -1165
rect -2109 -1199 -2093 -1165
rect -2035 -1199 -2019 -1165
rect -1851 -1199 -1835 -1165
rect -1777 -1199 -1761 -1165
rect -1593 -1199 -1577 -1165
rect -1519 -1199 -1503 -1165
rect -1335 -1199 -1319 -1165
rect -1261 -1199 -1245 -1165
rect -1077 -1199 -1061 -1165
rect -1003 -1199 -987 -1165
rect -819 -1199 -803 -1165
rect -745 -1199 -729 -1165
rect -561 -1199 -545 -1165
rect -487 -1199 -471 -1165
rect -303 -1199 -287 -1165
rect -229 -1199 -213 -1165
rect -45 -1199 -29 -1165
rect 29 -1199 45 -1165
rect 213 -1199 229 -1165
rect 287 -1199 303 -1165
rect 471 -1199 487 -1165
rect 545 -1199 561 -1165
rect 729 -1199 745 -1165
rect 803 -1199 819 -1165
rect 987 -1199 1003 -1165
rect 1061 -1199 1077 -1165
rect 1245 -1199 1261 -1165
rect 1319 -1199 1335 -1165
rect 1503 -1199 1519 -1165
rect 1577 -1199 1593 -1165
rect 1761 -1199 1777 -1165
rect 1835 -1199 1851 -1165
rect 2019 -1199 2035 -1165
rect 2093 -1199 2109 -1165
rect 2277 -1199 2293 -1165
rect 2351 -1199 2367 -1165
rect 2535 -1199 2551 -1165
rect 2609 -1199 2625 -1165
rect 2793 -1199 2809 -1165
rect 2867 -1199 2883 -1165
rect 3051 -1199 3067 -1165
rect 3125 -1199 3141 -1165
rect 3309 -1199 3325 -1165
rect 3383 -1199 3399 -1165
rect 3567 -1199 3583 -1165
rect -3583 -1307 -3567 -1273
rect -3399 -1307 -3383 -1273
rect -3325 -1307 -3309 -1273
rect -3141 -1307 -3125 -1273
rect -3067 -1307 -3051 -1273
rect -2883 -1307 -2867 -1273
rect -2809 -1307 -2793 -1273
rect -2625 -1307 -2609 -1273
rect -2551 -1307 -2535 -1273
rect -2367 -1307 -2351 -1273
rect -2293 -1307 -2277 -1273
rect -2109 -1307 -2093 -1273
rect -2035 -1307 -2019 -1273
rect -1851 -1307 -1835 -1273
rect -1777 -1307 -1761 -1273
rect -1593 -1307 -1577 -1273
rect -1519 -1307 -1503 -1273
rect -1335 -1307 -1319 -1273
rect -1261 -1307 -1245 -1273
rect -1077 -1307 -1061 -1273
rect -1003 -1307 -987 -1273
rect -819 -1307 -803 -1273
rect -745 -1307 -729 -1273
rect -561 -1307 -545 -1273
rect -487 -1307 -471 -1273
rect -303 -1307 -287 -1273
rect -229 -1307 -213 -1273
rect -45 -1307 -29 -1273
rect 29 -1307 45 -1273
rect 213 -1307 229 -1273
rect 287 -1307 303 -1273
rect 471 -1307 487 -1273
rect 545 -1307 561 -1273
rect 729 -1307 745 -1273
rect 803 -1307 819 -1273
rect 987 -1307 1003 -1273
rect 1061 -1307 1077 -1273
rect 1245 -1307 1261 -1273
rect 1319 -1307 1335 -1273
rect 1503 -1307 1519 -1273
rect 1577 -1307 1593 -1273
rect 1761 -1307 1777 -1273
rect 1835 -1307 1851 -1273
rect 2019 -1307 2035 -1273
rect 2093 -1307 2109 -1273
rect 2277 -1307 2293 -1273
rect 2351 -1307 2367 -1273
rect 2535 -1307 2551 -1273
rect 2609 -1307 2625 -1273
rect 2793 -1307 2809 -1273
rect 2867 -1307 2883 -1273
rect 3051 -1307 3067 -1273
rect 3125 -1307 3141 -1273
rect 3309 -1307 3325 -1273
rect 3383 -1307 3399 -1273
rect 3567 -1307 3583 -1273
rect -3629 -1366 -3595 -1350
rect -3629 -2358 -3595 -2342
rect -3371 -1366 -3337 -1350
rect -3371 -2358 -3337 -2342
rect -3113 -1366 -3079 -1350
rect -3113 -2358 -3079 -2342
rect -2855 -1366 -2821 -1350
rect -2855 -2358 -2821 -2342
rect -2597 -1366 -2563 -1350
rect -2597 -2358 -2563 -2342
rect -2339 -1366 -2305 -1350
rect -2339 -2358 -2305 -2342
rect -2081 -1366 -2047 -1350
rect -2081 -2358 -2047 -2342
rect -1823 -1366 -1789 -1350
rect -1823 -2358 -1789 -2342
rect -1565 -1366 -1531 -1350
rect -1565 -2358 -1531 -2342
rect -1307 -1366 -1273 -1350
rect -1307 -2358 -1273 -2342
rect -1049 -1366 -1015 -1350
rect -1049 -2358 -1015 -2342
rect -791 -1366 -757 -1350
rect -791 -2358 -757 -2342
rect -533 -1366 -499 -1350
rect -533 -2358 -499 -2342
rect -275 -1366 -241 -1350
rect -275 -2358 -241 -2342
rect -17 -1366 17 -1350
rect -17 -2358 17 -2342
rect 241 -1366 275 -1350
rect 241 -2358 275 -2342
rect 499 -1366 533 -1350
rect 499 -2358 533 -2342
rect 757 -1366 791 -1350
rect 757 -2358 791 -2342
rect 1015 -1366 1049 -1350
rect 1015 -2358 1049 -2342
rect 1273 -1366 1307 -1350
rect 1273 -2358 1307 -2342
rect 1531 -1366 1565 -1350
rect 1531 -2358 1565 -2342
rect 1789 -1366 1823 -1350
rect 1789 -2358 1823 -2342
rect 2047 -1366 2081 -1350
rect 2047 -2358 2081 -2342
rect 2305 -1366 2339 -1350
rect 2305 -2358 2339 -2342
rect 2563 -1366 2597 -1350
rect 2563 -2358 2597 -2342
rect 2821 -1366 2855 -1350
rect 2821 -2358 2855 -2342
rect 3079 -1366 3113 -1350
rect 3079 -2358 3113 -2342
rect 3337 -1366 3371 -1350
rect 3337 -2358 3371 -2342
rect 3595 -1366 3629 -1350
rect 3595 -2358 3629 -2342
rect -3583 -2435 -3567 -2401
rect -3399 -2435 -3383 -2401
rect -3325 -2435 -3309 -2401
rect -3141 -2435 -3125 -2401
rect -3067 -2435 -3051 -2401
rect -2883 -2435 -2867 -2401
rect -2809 -2435 -2793 -2401
rect -2625 -2435 -2609 -2401
rect -2551 -2435 -2535 -2401
rect -2367 -2435 -2351 -2401
rect -2293 -2435 -2277 -2401
rect -2109 -2435 -2093 -2401
rect -2035 -2435 -2019 -2401
rect -1851 -2435 -1835 -2401
rect -1777 -2435 -1761 -2401
rect -1593 -2435 -1577 -2401
rect -1519 -2435 -1503 -2401
rect -1335 -2435 -1319 -2401
rect -1261 -2435 -1245 -2401
rect -1077 -2435 -1061 -2401
rect -1003 -2435 -987 -2401
rect -819 -2435 -803 -2401
rect -745 -2435 -729 -2401
rect -561 -2435 -545 -2401
rect -487 -2435 -471 -2401
rect -303 -2435 -287 -2401
rect -229 -2435 -213 -2401
rect -45 -2435 -29 -2401
rect 29 -2435 45 -2401
rect 213 -2435 229 -2401
rect 287 -2435 303 -2401
rect 471 -2435 487 -2401
rect 545 -2435 561 -2401
rect 729 -2435 745 -2401
rect 803 -2435 819 -2401
rect 987 -2435 1003 -2401
rect 1061 -2435 1077 -2401
rect 1245 -2435 1261 -2401
rect 1319 -2435 1335 -2401
rect 1503 -2435 1519 -2401
rect 1577 -2435 1593 -2401
rect 1761 -2435 1777 -2401
rect 1835 -2435 1851 -2401
rect 2019 -2435 2035 -2401
rect 2093 -2435 2109 -2401
rect 2277 -2435 2293 -2401
rect 2351 -2435 2367 -2401
rect 2535 -2435 2551 -2401
rect 2609 -2435 2625 -2401
rect 2793 -2435 2809 -2401
rect 2867 -2435 2883 -2401
rect 3051 -2435 3067 -2401
rect 3125 -2435 3141 -2401
rect 3309 -2435 3325 -2401
rect 3383 -2435 3399 -2401
rect 3567 -2435 3583 -2401
rect -3763 -2539 -3729 -2477
rect 3729 -2539 3763 -2477
rect -3763 -2573 -3667 -2539
rect 3667 -2573 3763 -2539
<< viali >>
rect -3567 2401 -3399 2435
rect -3309 2401 -3141 2435
rect -3051 2401 -2883 2435
rect -2793 2401 -2625 2435
rect -2535 2401 -2367 2435
rect -2277 2401 -2109 2435
rect -2019 2401 -1851 2435
rect -1761 2401 -1593 2435
rect -1503 2401 -1335 2435
rect -1245 2401 -1077 2435
rect -987 2401 -819 2435
rect -729 2401 -561 2435
rect -471 2401 -303 2435
rect -213 2401 -45 2435
rect 45 2401 213 2435
rect 303 2401 471 2435
rect 561 2401 729 2435
rect 819 2401 987 2435
rect 1077 2401 1245 2435
rect 1335 2401 1503 2435
rect 1593 2401 1761 2435
rect 1851 2401 2019 2435
rect 2109 2401 2277 2435
rect 2367 2401 2535 2435
rect 2625 2401 2793 2435
rect 2883 2401 3051 2435
rect 3141 2401 3309 2435
rect 3399 2401 3567 2435
rect -3629 1366 -3595 2342
rect -3371 1366 -3337 2342
rect -3113 1366 -3079 2342
rect -2855 1366 -2821 2342
rect -2597 1366 -2563 2342
rect -2339 1366 -2305 2342
rect -2081 1366 -2047 2342
rect -1823 1366 -1789 2342
rect -1565 1366 -1531 2342
rect -1307 1366 -1273 2342
rect -1049 1366 -1015 2342
rect -791 1366 -757 2342
rect -533 1366 -499 2342
rect -275 1366 -241 2342
rect -17 1366 17 2342
rect 241 1366 275 2342
rect 499 1366 533 2342
rect 757 1366 791 2342
rect 1015 1366 1049 2342
rect 1273 1366 1307 2342
rect 1531 1366 1565 2342
rect 1789 1366 1823 2342
rect 2047 1366 2081 2342
rect 2305 1366 2339 2342
rect 2563 1366 2597 2342
rect 2821 1366 2855 2342
rect 3079 1366 3113 2342
rect 3337 1366 3371 2342
rect 3595 1366 3629 2342
rect -3567 1273 -3399 1307
rect -3309 1273 -3141 1307
rect -3051 1273 -2883 1307
rect -2793 1273 -2625 1307
rect -2535 1273 -2367 1307
rect -2277 1273 -2109 1307
rect -2019 1273 -1851 1307
rect -1761 1273 -1593 1307
rect -1503 1273 -1335 1307
rect -1245 1273 -1077 1307
rect -987 1273 -819 1307
rect -729 1273 -561 1307
rect -471 1273 -303 1307
rect -213 1273 -45 1307
rect 45 1273 213 1307
rect 303 1273 471 1307
rect 561 1273 729 1307
rect 819 1273 987 1307
rect 1077 1273 1245 1307
rect 1335 1273 1503 1307
rect 1593 1273 1761 1307
rect 1851 1273 2019 1307
rect 2109 1273 2277 1307
rect 2367 1273 2535 1307
rect 2625 1273 2793 1307
rect 2883 1273 3051 1307
rect 3141 1273 3309 1307
rect 3399 1273 3567 1307
rect -3567 1165 -3399 1199
rect -3309 1165 -3141 1199
rect -3051 1165 -2883 1199
rect -2793 1165 -2625 1199
rect -2535 1165 -2367 1199
rect -2277 1165 -2109 1199
rect -2019 1165 -1851 1199
rect -1761 1165 -1593 1199
rect -1503 1165 -1335 1199
rect -1245 1165 -1077 1199
rect -987 1165 -819 1199
rect -729 1165 -561 1199
rect -471 1165 -303 1199
rect -213 1165 -45 1199
rect 45 1165 213 1199
rect 303 1165 471 1199
rect 561 1165 729 1199
rect 819 1165 987 1199
rect 1077 1165 1245 1199
rect 1335 1165 1503 1199
rect 1593 1165 1761 1199
rect 1851 1165 2019 1199
rect 2109 1165 2277 1199
rect 2367 1165 2535 1199
rect 2625 1165 2793 1199
rect 2883 1165 3051 1199
rect 3141 1165 3309 1199
rect 3399 1165 3567 1199
rect -3629 130 -3595 1106
rect -3371 130 -3337 1106
rect -3113 130 -3079 1106
rect -2855 130 -2821 1106
rect -2597 130 -2563 1106
rect -2339 130 -2305 1106
rect -2081 130 -2047 1106
rect -1823 130 -1789 1106
rect -1565 130 -1531 1106
rect -1307 130 -1273 1106
rect -1049 130 -1015 1106
rect -791 130 -757 1106
rect -533 130 -499 1106
rect -275 130 -241 1106
rect -17 130 17 1106
rect 241 130 275 1106
rect 499 130 533 1106
rect 757 130 791 1106
rect 1015 130 1049 1106
rect 1273 130 1307 1106
rect 1531 130 1565 1106
rect 1789 130 1823 1106
rect 2047 130 2081 1106
rect 2305 130 2339 1106
rect 2563 130 2597 1106
rect 2821 130 2855 1106
rect 3079 130 3113 1106
rect 3337 130 3371 1106
rect 3595 130 3629 1106
rect -3567 37 -3399 71
rect -3309 37 -3141 71
rect -3051 37 -2883 71
rect -2793 37 -2625 71
rect -2535 37 -2367 71
rect -2277 37 -2109 71
rect -2019 37 -1851 71
rect -1761 37 -1593 71
rect -1503 37 -1335 71
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect 1335 37 1503 71
rect 1593 37 1761 71
rect 1851 37 2019 71
rect 2109 37 2277 71
rect 2367 37 2535 71
rect 2625 37 2793 71
rect 2883 37 3051 71
rect 3141 37 3309 71
rect 3399 37 3567 71
rect -3567 -71 -3399 -37
rect -3309 -71 -3141 -37
rect -3051 -71 -2883 -37
rect -2793 -71 -2625 -37
rect -2535 -71 -2367 -37
rect -2277 -71 -2109 -37
rect -2019 -71 -1851 -37
rect -1761 -71 -1593 -37
rect -1503 -71 -1335 -37
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect 1335 -71 1503 -37
rect 1593 -71 1761 -37
rect 1851 -71 2019 -37
rect 2109 -71 2277 -37
rect 2367 -71 2535 -37
rect 2625 -71 2793 -37
rect 2883 -71 3051 -37
rect 3141 -71 3309 -37
rect 3399 -71 3567 -37
rect -3629 -1106 -3595 -130
rect -3371 -1106 -3337 -130
rect -3113 -1106 -3079 -130
rect -2855 -1106 -2821 -130
rect -2597 -1106 -2563 -130
rect -2339 -1106 -2305 -130
rect -2081 -1106 -2047 -130
rect -1823 -1106 -1789 -130
rect -1565 -1106 -1531 -130
rect -1307 -1106 -1273 -130
rect -1049 -1106 -1015 -130
rect -791 -1106 -757 -130
rect -533 -1106 -499 -130
rect -275 -1106 -241 -130
rect -17 -1106 17 -130
rect 241 -1106 275 -130
rect 499 -1106 533 -130
rect 757 -1106 791 -130
rect 1015 -1106 1049 -130
rect 1273 -1106 1307 -130
rect 1531 -1106 1565 -130
rect 1789 -1106 1823 -130
rect 2047 -1106 2081 -130
rect 2305 -1106 2339 -130
rect 2563 -1106 2597 -130
rect 2821 -1106 2855 -130
rect 3079 -1106 3113 -130
rect 3337 -1106 3371 -130
rect 3595 -1106 3629 -130
rect -3567 -1199 -3399 -1165
rect -3309 -1199 -3141 -1165
rect -3051 -1199 -2883 -1165
rect -2793 -1199 -2625 -1165
rect -2535 -1199 -2367 -1165
rect -2277 -1199 -2109 -1165
rect -2019 -1199 -1851 -1165
rect -1761 -1199 -1593 -1165
rect -1503 -1199 -1335 -1165
rect -1245 -1199 -1077 -1165
rect -987 -1199 -819 -1165
rect -729 -1199 -561 -1165
rect -471 -1199 -303 -1165
rect -213 -1199 -45 -1165
rect 45 -1199 213 -1165
rect 303 -1199 471 -1165
rect 561 -1199 729 -1165
rect 819 -1199 987 -1165
rect 1077 -1199 1245 -1165
rect 1335 -1199 1503 -1165
rect 1593 -1199 1761 -1165
rect 1851 -1199 2019 -1165
rect 2109 -1199 2277 -1165
rect 2367 -1199 2535 -1165
rect 2625 -1199 2793 -1165
rect 2883 -1199 3051 -1165
rect 3141 -1199 3309 -1165
rect 3399 -1199 3567 -1165
rect -3567 -1307 -3399 -1273
rect -3309 -1307 -3141 -1273
rect -3051 -1307 -2883 -1273
rect -2793 -1307 -2625 -1273
rect -2535 -1307 -2367 -1273
rect -2277 -1307 -2109 -1273
rect -2019 -1307 -1851 -1273
rect -1761 -1307 -1593 -1273
rect -1503 -1307 -1335 -1273
rect -1245 -1307 -1077 -1273
rect -987 -1307 -819 -1273
rect -729 -1307 -561 -1273
rect -471 -1307 -303 -1273
rect -213 -1307 -45 -1273
rect 45 -1307 213 -1273
rect 303 -1307 471 -1273
rect 561 -1307 729 -1273
rect 819 -1307 987 -1273
rect 1077 -1307 1245 -1273
rect 1335 -1307 1503 -1273
rect 1593 -1307 1761 -1273
rect 1851 -1307 2019 -1273
rect 2109 -1307 2277 -1273
rect 2367 -1307 2535 -1273
rect 2625 -1307 2793 -1273
rect 2883 -1307 3051 -1273
rect 3141 -1307 3309 -1273
rect 3399 -1307 3567 -1273
rect -3629 -2342 -3595 -1366
rect -3371 -2342 -3337 -1366
rect -3113 -2342 -3079 -1366
rect -2855 -2342 -2821 -1366
rect -2597 -2342 -2563 -1366
rect -2339 -2342 -2305 -1366
rect -2081 -2342 -2047 -1366
rect -1823 -2342 -1789 -1366
rect -1565 -2342 -1531 -1366
rect -1307 -2342 -1273 -1366
rect -1049 -2342 -1015 -1366
rect -791 -2342 -757 -1366
rect -533 -2342 -499 -1366
rect -275 -2342 -241 -1366
rect -17 -2342 17 -1366
rect 241 -2342 275 -1366
rect 499 -2342 533 -1366
rect 757 -2342 791 -1366
rect 1015 -2342 1049 -1366
rect 1273 -2342 1307 -1366
rect 1531 -2342 1565 -1366
rect 1789 -2342 1823 -1366
rect 2047 -2342 2081 -1366
rect 2305 -2342 2339 -1366
rect 2563 -2342 2597 -1366
rect 2821 -2342 2855 -1366
rect 3079 -2342 3113 -1366
rect 3337 -2342 3371 -1366
rect 3595 -2342 3629 -1366
rect -3567 -2435 -3399 -2401
rect -3309 -2435 -3141 -2401
rect -3051 -2435 -2883 -2401
rect -2793 -2435 -2625 -2401
rect -2535 -2435 -2367 -2401
rect -2277 -2435 -2109 -2401
rect -2019 -2435 -1851 -2401
rect -1761 -2435 -1593 -2401
rect -1503 -2435 -1335 -2401
rect -1245 -2435 -1077 -2401
rect -987 -2435 -819 -2401
rect -729 -2435 -561 -2401
rect -471 -2435 -303 -2401
rect -213 -2435 -45 -2401
rect 45 -2435 213 -2401
rect 303 -2435 471 -2401
rect 561 -2435 729 -2401
rect 819 -2435 987 -2401
rect 1077 -2435 1245 -2401
rect 1335 -2435 1503 -2401
rect 1593 -2435 1761 -2401
rect 1851 -2435 2019 -2401
rect 2109 -2435 2277 -2401
rect 2367 -2435 2535 -2401
rect 2625 -2435 2793 -2401
rect 2883 -2435 3051 -2401
rect 3141 -2435 3309 -2401
rect 3399 -2435 3567 -2401
<< metal1 >>
rect -3579 2435 -3387 2441
rect -3579 2401 -3567 2435
rect -3399 2401 -3387 2435
rect -3579 2395 -3387 2401
rect -3321 2435 -3129 2441
rect -3321 2401 -3309 2435
rect -3141 2401 -3129 2435
rect -3321 2395 -3129 2401
rect -3063 2435 -2871 2441
rect -3063 2401 -3051 2435
rect -2883 2401 -2871 2435
rect -3063 2395 -2871 2401
rect -2805 2435 -2613 2441
rect -2805 2401 -2793 2435
rect -2625 2401 -2613 2435
rect -2805 2395 -2613 2401
rect -2547 2435 -2355 2441
rect -2547 2401 -2535 2435
rect -2367 2401 -2355 2435
rect -2547 2395 -2355 2401
rect -2289 2435 -2097 2441
rect -2289 2401 -2277 2435
rect -2109 2401 -2097 2435
rect -2289 2395 -2097 2401
rect -2031 2435 -1839 2441
rect -2031 2401 -2019 2435
rect -1851 2401 -1839 2435
rect -2031 2395 -1839 2401
rect -1773 2435 -1581 2441
rect -1773 2401 -1761 2435
rect -1593 2401 -1581 2435
rect -1773 2395 -1581 2401
rect -1515 2435 -1323 2441
rect -1515 2401 -1503 2435
rect -1335 2401 -1323 2435
rect -1515 2395 -1323 2401
rect -1257 2435 -1065 2441
rect -1257 2401 -1245 2435
rect -1077 2401 -1065 2435
rect -1257 2395 -1065 2401
rect -999 2435 -807 2441
rect -999 2401 -987 2435
rect -819 2401 -807 2435
rect -999 2395 -807 2401
rect -741 2435 -549 2441
rect -741 2401 -729 2435
rect -561 2401 -549 2435
rect -741 2395 -549 2401
rect -483 2435 -291 2441
rect -483 2401 -471 2435
rect -303 2401 -291 2435
rect -483 2395 -291 2401
rect -225 2435 -33 2441
rect -225 2401 -213 2435
rect -45 2401 -33 2435
rect -225 2395 -33 2401
rect 33 2435 225 2441
rect 33 2401 45 2435
rect 213 2401 225 2435
rect 33 2395 225 2401
rect 291 2435 483 2441
rect 291 2401 303 2435
rect 471 2401 483 2435
rect 291 2395 483 2401
rect 549 2435 741 2441
rect 549 2401 561 2435
rect 729 2401 741 2435
rect 549 2395 741 2401
rect 807 2435 999 2441
rect 807 2401 819 2435
rect 987 2401 999 2435
rect 807 2395 999 2401
rect 1065 2435 1257 2441
rect 1065 2401 1077 2435
rect 1245 2401 1257 2435
rect 1065 2395 1257 2401
rect 1323 2435 1515 2441
rect 1323 2401 1335 2435
rect 1503 2401 1515 2435
rect 1323 2395 1515 2401
rect 1581 2435 1773 2441
rect 1581 2401 1593 2435
rect 1761 2401 1773 2435
rect 1581 2395 1773 2401
rect 1839 2435 2031 2441
rect 1839 2401 1851 2435
rect 2019 2401 2031 2435
rect 1839 2395 2031 2401
rect 2097 2435 2289 2441
rect 2097 2401 2109 2435
rect 2277 2401 2289 2435
rect 2097 2395 2289 2401
rect 2355 2435 2547 2441
rect 2355 2401 2367 2435
rect 2535 2401 2547 2435
rect 2355 2395 2547 2401
rect 2613 2435 2805 2441
rect 2613 2401 2625 2435
rect 2793 2401 2805 2435
rect 2613 2395 2805 2401
rect 2871 2435 3063 2441
rect 2871 2401 2883 2435
rect 3051 2401 3063 2435
rect 2871 2395 3063 2401
rect 3129 2435 3321 2441
rect 3129 2401 3141 2435
rect 3309 2401 3321 2435
rect 3129 2395 3321 2401
rect 3387 2435 3579 2441
rect 3387 2401 3399 2435
rect 3567 2401 3579 2435
rect 3387 2395 3579 2401
rect -3635 2342 -3589 2354
rect -3635 1366 -3629 2342
rect -3595 1366 -3589 2342
rect -3635 1354 -3589 1366
rect -3377 2342 -3331 2354
rect -3377 1366 -3371 2342
rect -3337 1366 -3331 2342
rect -3377 1354 -3331 1366
rect -3119 2342 -3073 2354
rect -3119 1366 -3113 2342
rect -3079 1366 -3073 2342
rect -3119 1354 -3073 1366
rect -2861 2342 -2815 2354
rect -2861 1366 -2855 2342
rect -2821 1366 -2815 2342
rect -2861 1354 -2815 1366
rect -2603 2342 -2557 2354
rect -2603 1366 -2597 2342
rect -2563 1366 -2557 2342
rect -2603 1354 -2557 1366
rect -2345 2342 -2299 2354
rect -2345 1366 -2339 2342
rect -2305 1366 -2299 2342
rect -2345 1354 -2299 1366
rect -2087 2342 -2041 2354
rect -2087 1366 -2081 2342
rect -2047 1366 -2041 2342
rect -2087 1354 -2041 1366
rect -1829 2342 -1783 2354
rect -1829 1366 -1823 2342
rect -1789 1366 -1783 2342
rect -1829 1354 -1783 1366
rect -1571 2342 -1525 2354
rect -1571 1366 -1565 2342
rect -1531 1366 -1525 2342
rect -1571 1354 -1525 1366
rect -1313 2342 -1267 2354
rect -1313 1366 -1307 2342
rect -1273 1366 -1267 2342
rect -1313 1354 -1267 1366
rect -1055 2342 -1009 2354
rect -1055 1366 -1049 2342
rect -1015 1366 -1009 2342
rect -1055 1354 -1009 1366
rect -797 2342 -751 2354
rect -797 1366 -791 2342
rect -757 1366 -751 2342
rect -797 1354 -751 1366
rect -539 2342 -493 2354
rect -539 1366 -533 2342
rect -499 1366 -493 2342
rect -539 1354 -493 1366
rect -281 2342 -235 2354
rect -281 1366 -275 2342
rect -241 1366 -235 2342
rect -281 1354 -235 1366
rect -23 2342 23 2354
rect -23 1366 -17 2342
rect 17 1366 23 2342
rect -23 1354 23 1366
rect 235 2342 281 2354
rect 235 1366 241 2342
rect 275 1366 281 2342
rect 235 1354 281 1366
rect 493 2342 539 2354
rect 493 1366 499 2342
rect 533 1366 539 2342
rect 493 1354 539 1366
rect 751 2342 797 2354
rect 751 1366 757 2342
rect 791 1366 797 2342
rect 751 1354 797 1366
rect 1009 2342 1055 2354
rect 1009 1366 1015 2342
rect 1049 1366 1055 2342
rect 1009 1354 1055 1366
rect 1267 2342 1313 2354
rect 1267 1366 1273 2342
rect 1307 1366 1313 2342
rect 1267 1354 1313 1366
rect 1525 2342 1571 2354
rect 1525 1366 1531 2342
rect 1565 1366 1571 2342
rect 1525 1354 1571 1366
rect 1783 2342 1829 2354
rect 1783 1366 1789 2342
rect 1823 1366 1829 2342
rect 1783 1354 1829 1366
rect 2041 2342 2087 2354
rect 2041 1366 2047 2342
rect 2081 1366 2087 2342
rect 2041 1354 2087 1366
rect 2299 2342 2345 2354
rect 2299 1366 2305 2342
rect 2339 1366 2345 2342
rect 2299 1354 2345 1366
rect 2557 2342 2603 2354
rect 2557 1366 2563 2342
rect 2597 1366 2603 2342
rect 2557 1354 2603 1366
rect 2815 2342 2861 2354
rect 2815 1366 2821 2342
rect 2855 1366 2861 2342
rect 2815 1354 2861 1366
rect 3073 2342 3119 2354
rect 3073 1366 3079 2342
rect 3113 1366 3119 2342
rect 3073 1354 3119 1366
rect 3331 2342 3377 2354
rect 3331 1366 3337 2342
rect 3371 1366 3377 2342
rect 3331 1354 3377 1366
rect 3589 2342 3635 2354
rect 3589 1366 3595 2342
rect 3629 1366 3635 2342
rect 3589 1354 3635 1366
rect -3579 1307 -3387 1313
rect -3579 1273 -3567 1307
rect -3399 1273 -3387 1307
rect -3579 1267 -3387 1273
rect -3321 1307 -3129 1313
rect -3321 1273 -3309 1307
rect -3141 1273 -3129 1307
rect -3321 1267 -3129 1273
rect -3063 1307 -2871 1313
rect -3063 1273 -3051 1307
rect -2883 1273 -2871 1307
rect -3063 1267 -2871 1273
rect -2805 1307 -2613 1313
rect -2805 1273 -2793 1307
rect -2625 1273 -2613 1307
rect -2805 1267 -2613 1273
rect -2547 1307 -2355 1313
rect -2547 1273 -2535 1307
rect -2367 1273 -2355 1307
rect -2547 1267 -2355 1273
rect -2289 1307 -2097 1313
rect -2289 1273 -2277 1307
rect -2109 1273 -2097 1307
rect -2289 1267 -2097 1273
rect -2031 1307 -1839 1313
rect -2031 1273 -2019 1307
rect -1851 1273 -1839 1307
rect -2031 1267 -1839 1273
rect -1773 1307 -1581 1313
rect -1773 1273 -1761 1307
rect -1593 1273 -1581 1307
rect -1773 1267 -1581 1273
rect -1515 1307 -1323 1313
rect -1515 1273 -1503 1307
rect -1335 1273 -1323 1307
rect -1515 1267 -1323 1273
rect -1257 1307 -1065 1313
rect -1257 1273 -1245 1307
rect -1077 1273 -1065 1307
rect -1257 1267 -1065 1273
rect -999 1307 -807 1313
rect -999 1273 -987 1307
rect -819 1273 -807 1307
rect -999 1267 -807 1273
rect -741 1307 -549 1313
rect -741 1273 -729 1307
rect -561 1273 -549 1307
rect -741 1267 -549 1273
rect -483 1307 -291 1313
rect -483 1273 -471 1307
rect -303 1273 -291 1307
rect -483 1267 -291 1273
rect -225 1307 -33 1313
rect -225 1273 -213 1307
rect -45 1273 -33 1307
rect -225 1267 -33 1273
rect 33 1307 225 1313
rect 33 1273 45 1307
rect 213 1273 225 1307
rect 33 1267 225 1273
rect 291 1307 483 1313
rect 291 1273 303 1307
rect 471 1273 483 1307
rect 291 1267 483 1273
rect 549 1307 741 1313
rect 549 1273 561 1307
rect 729 1273 741 1307
rect 549 1267 741 1273
rect 807 1307 999 1313
rect 807 1273 819 1307
rect 987 1273 999 1307
rect 807 1267 999 1273
rect 1065 1307 1257 1313
rect 1065 1273 1077 1307
rect 1245 1273 1257 1307
rect 1065 1267 1257 1273
rect 1323 1307 1515 1313
rect 1323 1273 1335 1307
rect 1503 1273 1515 1307
rect 1323 1267 1515 1273
rect 1581 1307 1773 1313
rect 1581 1273 1593 1307
rect 1761 1273 1773 1307
rect 1581 1267 1773 1273
rect 1839 1307 2031 1313
rect 1839 1273 1851 1307
rect 2019 1273 2031 1307
rect 1839 1267 2031 1273
rect 2097 1307 2289 1313
rect 2097 1273 2109 1307
rect 2277 1273 2289 1307
rect 2097 1267 2289 1273
rect 2355 1307 2547 1313
rect 2355 1273 2367 1307
rect 2535 1273 2547 1307
rect 2355 1267 2547 1273
rect 2613 1307 2805 1313
rect 2613 1273 2625 1307
rect 2793 1273 2805 1307
rect 2613 1267 2805 1273
rect 2871 1307 3063 1313
rect 2871 1273 2883 1307
rect 3051 1273 3063 1307
rect 2871 1267 3063 1273
rect 3129 1307 3321 1313
rect 3129 1273 3141 1307
rect 3309 1273 3321 1307
rect 3129 1267 3321 1273
rect 3387 1307 3579 1313
rect 3387 1273 3399 1307
rect 3567 1273 3579 1307
rect 3387 1267 3579 1273
rect -3579 1199 -3387 1205
rect -3579 1165 -3567 1199
rect -3399 1165 -3387 1199
rect -3579 1159 -3387 1165
rect -3321 1199 -3129 1205
rect -3321 1165 -3309 1199
rect -3141 1165 -3129 1199
rect -3321 1159 -3129 1165
rect -3063 1199 -2871 1205
rect -3063 1165 -3051 1199
rect -2883 1165 -2871 1199
rect -3063 1159 -2871 1165
rect -2805 1199 -2613 1205
rect -2805 1165 -2793 1199
rect -2625 1165 -2613 1199
rect -2805 1159 -2613 1165
rect -2547 1199 -2355 1205
rect -2547 1165 -2535 1199
rect -2367 1165 -2355 1199
rect -2547 1159 -2355 1165
rect -2289 1199 -2097 1205
rect -2289 1165 -2277 1199
rect -2109 1165 -2097 1199
rect -2289 1159 -2097 1165
rect -2031 1199 -1839 1205
rect -2031 1165 -2019 1199
rect -1851 1165 -1839 1199
rect -2031 1159 -1839 1165
rect -1773 1199 -1581 1205
rect -1773 1165 -1761 1199
rect -1593 1165 -1581 1199
rect -1773 1159 -1581 1165
rect -1515 1199 -1323 1205
rect -1515 1165 -1503 1199
rect -1335 1165 -1323 1199
rect -1515 1159 -1323 1165
rect -1257 1199 -1065 1205
rect -1257 1165 -1245 1199
rect -1077 1165 -1065 1199
rect -1257 1159 -1065 1165
rect -999 1199 -807 1205
rect -999 1165 -987 1199
rect -819 1165 -807 1199
rect -999 1159 -807 1165
rect -741 1199 -549 1205
rect -741 1165 -729 1199
rect -561 1165 -549 1199
rect -741 1159 -549 1165
rect -483 1199 -291 1205
rect -483 1165 -471 1199
rect -303 1165 -291 1199
rect -483 1159 -291 1165
rect -225 1199 -33 1205
rect -225 1165 -213 1199
rect -45 1165 -33 1199
rect -225 1159 -33 1165
rect 33 1199 225 1205
rect 33 1165 45 1199
rect 213 1165 225 1199
rect 33 1159 225 1165
rect 291 1199 483 1205
rect 291 1165 303 1199
rect 471 1165 483 1199
rect 291 1159 483 1165
rect 549 1199 741 1205
rect 549 1165 561 1199
rect 729 1165 741 1199
rect 549 1159 741 1165
rect 807 1199 999 1205
rect 807 1165 819 1199
rect 987 1165 999 1199
rect 807 1159 999 1165
rect 1065 1199 1257 1205
rect 1065 1165 1077 1199
rect 1245 1165 1257 1199
rect 1065 1159 1257 1165
rect 1323 1199 1515 1205
rect 1323 1165 1335 1199
rect 1503 1165 1515 1199
rect 1323 1159 1515 1165
rect 1581 1199 1773 1205
rect 1581 1165 1593 1199
rect 1761 1165 1773 1199
rect 1581 1159 1773 1165
rect 1839 1199 2031 1205
rect 1839 1165 1851 1199
rect 2019 1165 2031 1199
rect 1839 1159 2031 1165
rect 2097 1199 2289 1205
rect 2097 1165 2109 1199
rect 2277 1165 2289 1199
rect 2097 1159 2289 1165
rect 2355 1199 2547 1205
rect 2355 1165 2367 1199
rect 2535 1165 2547 1199
rect 2355 1159 2547 1165
rect 2613 1199 2805 1205
rect 2613 1165 2625 1199
rect 2793 1165 2805 1199
rect 2613 1159 2805 1165
rect 2871 1199 3063 1205
rect 2871 1165 2883 1199
rect 3051 1165 3063 1199
rect 2871 1159 3063 1165
rect 3129 1199 3321 1205
rect 3129 1165 3141 1199
rect 3309 1165 3321 1199
rect 3129 1159 3321 1165
rect 3387 1199 3579 1205
rect 3387 1165 3399 1199
rect 3567 1165 3579 1199
rect 3387 1159 3579 1165
rect -3635 1106 -3589 1118
rect -3635 130 -3629 1106
rect -3595 130 -3589 1106
rect -3635 118 -3589 130
rect -3377 1106 -3331 1118
rect -3377 130 -3371 1106
rect -3337 130 -3331 1106
rect -3377 118 -3331 130
rect -3119 1106 -3073 1118
rect -3119 130 -3113 1106
rect -3079 130 -3073 1106
rect -3119 118 -3073 130
rect -2861 1106 -2815 1118
rect -2861 130 -2855 1106
rect -2821 130 -2815 1106
rect -2861 118 -2815 130
rect -2603 1106 -2557 1118
rect -2603 130 -2597 1106
rect -2563 130 -2557 1106
rect -2603 118 -2557 130
rect -2345 1106 -2299 1118
rect -2345 130 -2339 1106
rect -2305 130 -2299 1106
rect -2345 118 -2299 130
rect -2087 1106 -2041 1118
rect -2087 130 -2081 1106
rect -2047 130 -2041 1106
rect -2087 118 -2041 130
rect -1829 1106 -1783 1118
rect -1829 130 -1823 1106
rect -1789 130 -1783 1106
rect -1829 118 -1783 130
rect -1571 1106 -1525 1118
rect -1571 130 -1565 1106
rect -1531 130 -1525 1106
rect -1571 118 -1525 130
rect -1313 1106 -1267 1118
rect -1313 130 -1307 1106
rect -1273 130 -1267 1106
rect -1313 118 -1267 130
rect -1055 1106 -1009 1118
rect -1055 130 -1049 1106
rect -1015 130 -1009 1106
rect -1055 118 -1009 130
rect -797 1106 -751 1118
rect -797 130 -791 1106
rect -757 130 -751 1106
rect -797 118 -751 130
rect -539 1106 -493 1118
rect -539 130 -533 1106
rect -499 130 -493 1106
rect -539 118 -493 130
rect -281 1106 -235 1118
rect -281 130 -275 1106
rect -241 130 -235 1106
rect -281 118 -235 130
rect -23 1106 23 1118
rect -23 130 -17 1106
rect 17 130 23 1106
rect -23 118 23 130
rect 235 1106 281 1118
rect 235 130 241 1106
rect 275 130 281 1106
rect 235 118 281 130
rect 493 1106 539 1118
rect 493 130 499 1106
rect 533 130 539 1106
rect 493 118 539 130
rect 751 1106 797 1118
rect 751 130 757 1106
rect 791 130 797 1106
rect 751 118 797 130
rect 1009 1106 1055 1118
rect 1009 130 1015 1106
rect 1049 130 1055 1106
rect 1009 118 1055 130
rect 1267 1106 1313 1118
rect 1267 130 1273 1106
rect 1307 130 1313 1106
rect 1267 118 1313 130
rect 1525 1106 1571 1118
rect 1525 130 1531 1106
rect 1565 130 1571 1106
rect 1525 118 1571 130
rect 1783 1106 1829 1118
rect 1783 130 1789 1106
rect 1823 130 1829 1106
rect 1783 118 1829 130
rect 2041 1106 2087 1118
rect 2041 130 2047 1106
rect 2081 130 2087 1106
rect 2041 118 2087 130
rect 2299 1106 2345 1118
rect 2299 130 2305 1106
rect 2339 130 2345 1106
rect 2299 118 2345 130
rect 2557 1106 2603 1118
rect 2557 130 2563 1106
rect 2597 130 2603 1106
rect 2557 118 2603 130
rect 2815 1106 2861 1118
rect 2815 130 2821 1106
rect 2855 130 2861 1106
rect 2815 118 2861 130
rect 3073 1106 3119 1118
rect 3073 130 3079 1106
rect 3113 130 3119 1106
rect 3073 118 3119 130
rect 3331 1106 3377 1118
rect 3331 130 3337 1106
rect 3371 130 3377 1106
rect 3331 118 3377 130
rect 3589 1106 3635 1118
rect 3589 130 3595 1106
rect 3629 130 3635 1106
rect 3589 118 3635 130
rect -3579 71 -3387 77
rect -3579 37 -3567 71
rect -3399 37 -3387 71
rect -3579 31 -3387 37
rect -3321 71 -3129 77
rect -3321 37 -3309 71
rect -3141 37 -3129 71
rect -3321 31 -3129 37
rect -3063 71 -2871 77
rect -3063 37 -3051 71
rect -2883 37 -2871 71
rect -3063 31 -2871 37
rect -2805 71 -2613 77
rect -2805 37 -2793 71
rect -2625 37 -2613 71
rect -2805 31 -2613 37
rect -2547 71 -2355 77
rect -2547 37 -2535 71
rect -2367 37 -2355 71
rect -2547 31 -2355 37
rect -2289 71 -2097 77
rect -2289 37 -2277 71
rect -2109 37 -2097 71
rect -2289 31 -2097 37
rect -2031 71 -1839 77
rect -2031 37 -2019 71
rect -1851 37 -1839 71
rect -2031 31 -1839 37
rect -1773 71 -1581 77
rect -1773 37 -1761 71
rect -1593 37 -1581 71
rect -1773 31 -1581 37
rect -1515 71 -1323 77
rect -1515 37 -1503 71
rect -1335 37 -1323 71
rect -1515 31 -1323 37
rect -1257 71 -1065 77
rect -1257 37 -1245 71
rect -1077 37 -1065 71
rect -1257 31 -1065 37
rect -999 71 -807 77
rect -999 37 -987 71
rect -819 37 -807 71
rect -999 31 -807 37
rect -741 71 -549 77
rect -741 37 -729 71
rect -561 37 -549 71
rect -741 31 -549 37
rect -483 71 -291 77
rect -483 37 -471 71
rect -303 37 -291 71
rect -483 31 -291 37
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect 291 71 483 77
rect 291 37 303 71
rect 471 37 483 71
rect 291 31 483 37
rect 549 71 741 77
rect 549 37 561 71
rect 729 37 741 71
rect 549 31 741 37
rect 807 71 999 77
rect 807 37 819 71
rect 987 37 999 71
rect 807 31 999 37
rect 1065 71 1257 77
rect 1065 37 1077 71
rect 1245 37 1257 71
rect 1065 31 1257 37
rect 1323 71 1515 77
rect 1323 37 1335 71
rect 1503 37 1515 71
rect 1323 31 1515 37
rect 1581 71 1773 77
rect 1581 37 1593 71
rect 1761 37 1773 71
rect 1581 31 1773 37
rect 1839 71 2031 77
rect 1839 37 1851 71
rect 2019 37 2031 71
rect 1839 31 2031 37
rect 2097 71 2289 77
rect 2097 37 2109 71
rect 2277 37 2289 71
rect 2097 31 2289 37
rect 2355 71 2547 77
rect 2355 37 2367 71
rect 2535 37 2547 71
rect 2355 31 2547 37
rect 2613 71 2805 77
rect 2613 37 2625 71
rect 2793 37 2805 71
rect 2613 31 2805 37
rect 2871 71 3063 77
rect 2871 37 2883 71
rect 3051 37 3063 71
rect 2871 31 3063 37
rect 3129 71 3321 77
rect 3129 37 3141 71
rect 3309 37 3321 71
rect 3129 31 3321 37
rect 3387 71 3579 77
rect 3387 37 3399 71
rect 3567 37 3579 71
rect 3387 31 3579 37
rect -3579 -37 -3387 -31
rect -3579 -71 -3567 -37
rect -3399 -71 -3387 -37
rect -3579 -77 -3387 -71
rect -3321 -37 -3129 -31
rect -3321 -71 -3309 -37
rect -3141 -71 -3129 -37
rect -3321 -77 -3129 -71
rect -3063 -37 -2871 -31
rect -3063 -71 -3051 -37
rect -2883 -71 -2871 -37
rect -3063 -77 -2871 -71
rect -2805 -37 -2613 -31
rect -2805 -71 -2793 -37
rect -2625 -71 -2613 -37
rect -2805 -77 -2613 -71
rect -2547 -37 -2355 -31
rect -2547 -71 -2535 -37
rect -2367 -71 -2355 -37
rect -2547 -77 -2355 -71
rect -2289 -37 -2097 -31
rect -2289 -71 -2277 -37
rect -2109 -71 -2097 -37
rect -2289 -77 -2097 -71
rect -2031 -37 -1839 -31
rect -2031 -71 -2019 -37
rect -1851 -71 -1839 -37
rect -2031 -77 -1839 -71
rect -1773 -37 -1581 -31
rect -1773 -71 -1761 -37
rect -1593 -71 -1581 -37
rect -1773 -77 -1581 -71
rect -1515 -37 -1323 -31
rect -1515 -71 -1503 -37
rect -1335 -71 -1323 -37
rect -1515 -77 -1323 -71
rect -1257 -37 -1065 -31
rect -1257 -71 -1245 -37
rect -1077 -71 -1065 -37
rect -1257 -77 -1065 -71
rect -999 -37 -807 -31
rect -999 -71 -987 -37
rect -819 -71 -807 -37
rect -999 -77 -807 -71
rect -741 -37 -549 -31
rect -741 -71 -729 -37
rect -561 -71 -549 -37
rect -741 -77 -549 -71
rect -483 -37 -291 -31
rect -483 -71 -471 -37
rect -303 -71 -291 -37
rect -483 -77 -291 -71
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect 291 -37 483 -31
rect 291 -71 303 -37
rect 471 -71 483 -37
rect 291 -77 483 -71
rect 549 -37 741 -31
rect 549 -71 561 -37
rect 729 -71 741 -37
rect 549 -77 741 -71
rect 807 -37 999 -31
rect 807 -71 819 -37
rect 987 -71 999 -37
rect 807 -77 999 -71
rect 1065 -37 1257 -31
rect 1065 -71 1077 -37
rect 1245 -71 1257 -37
rect 1065 -77 1257 -71
rect 1323 -37 1515 -31
rect 1323 -71 1335 -37
rect 1503 -71 1515 -37
rect 1323 -77 1515 -71
rect 1581 -37 1773 -31
rect 1581 -71 1593 -37
rect 1761 -71 1773 -37
rect 1581 -77 1773 -71
rect 1839 -37 2031 -31
rect 1839 -71 1851 -37
rect 2019 -71 2031 -37
rect 1839 -77 2031 -71
rect 2097 -37 2289 -31
rect 2097 -71 2109 -37
rect 2277 -71 2289 -37
rect 2097 -77 2289 -71
rect 2355 -37 2547 -31
rect 2355 -71 2367 -37
rect 2535 -71 2547 -37
rect 2355 -77 2547 -71
rect 2613 -37 2805 -31
rect 2613 -71 2625 -37
rect 2793 -71 2805 -37
rect 2613 -77 2805 -71
rect 2871 -37 3063 -31
rect 2871 -71 2883 -37
rect 3051 -71 3063 -37
rect 2871 -77 3063 -71
rect 3129 -37 3321 -31
rect 3129 -71 3141 -37
rect 3309 -71 3321 -37
rect 3129 -77 3321 -71
rect 3387 -37 3579 -31
rect 3387 -71 3399 -37
rect 3567 -71 3579 -37
rect 3387 -77 3579 -71
rect -3635 -130 -3589 -118
rect -3635 -1106 -3629 -130
rect -3595 -1106 -3589 -130
rect -3635 -1118 -3589 -1106
rect -3377 -130 -3331 -118
rect -3377 -1106 -3371 -130
rect -3337 -1106 -3331 -130
rect -3377 -1118 -3331 -1106
rect -3119 -130 -3073 -118
rect -3119 -1106 -3113 -130
rect -3079 -1106 -3073 -130
rect -3119 -1118 -3073 -1106
rect -2861 -130 -2815 -118
rect -2861 -1106 -2855 -130
rect -2821 -1106 -2815 -130
rect -2861 -1118 -2815 -1106
rect -2603 -130 -2557 -118
rect -2603 -1106 -2597 -130
rect -2563 -1106 -2557 -130
rect -2603 -1118 -2557 -1106
rect -2345 -130 -2299 -118
rect -2345 -1106 -2339 -130
rect -2305 -1106 -2299 -130
rect -2345 -1118 -2299 -1106
rect -2087 -130 -2041 -118
rect -2087 -1106 -2081 -130
rect -2047 -1106 -2041 -130
rect -2087 -1118 -2041 -1106
rect -1829 -130 -1783 -118
rect -1829 -1106 -1823 -130
rect -1789 -1106 -1783 -130
rect -1829 -1118 -1783 -1106
rect -1571 -130 -1525 -118
rect -1571 -1106 -1565 -130
rect -1531 -1106 -1525 -130
rect -1571 -1118 -1525 -1106
rect -1313 -130 -1267 -118
rect -1313 -1106 -1307 -130
rect -1273 -1106 -1267 -130
rect -1313 -1118 -1267 -1106
rect -1055 -130 -1009 -118
rect -1055 -1106 -1049 -130
rect -1015 -1106 -1009 -130
rect -1055 -1118 -1009 -1106
rect -797 -130 -751 -118
rect -797 -1106 -791 -130
rect -757 -1106 -751 -130
rect -797 -1118 -751 -1106
rect -539 -130 -493 -118
rect -539 -1106 -533 -130
rect -499 -1106 -493 -130
rect -539 -1118 -493 -1106
rect -281 -130 -235 -118
rect -281 -1106 -275 -130
rect -241 -1106 -235 -130
rect -281 -1118 -235 -1106
rect -23 -130 23 -118
rect -23 -1106 -17 -130
rect 17 -1106 23 -130
rect -23 -1118 23 -1106
rect 235 -130 281 -118
rect 235 -1106 241 -130
rect 275 -1106 281 -130
rect 235 -1118 281 -1106
rect 493 -130 539 -118
rect 493 -1106 499 -130
rect 533 -1106 539 -130
rect 493 -1118 539 -1106
rect 751 -130 797 -118
rect 751 -1106 757 -130
rect 791 -1106 797 -130
rect 751 -1118 797 -1106
rect 1009 -130 1055 -118
rect 1009 -1106 1015 -130
rect 1049 -1106 1055 -130
rect 1009 -1118 1055 -1106
rect 1267 -130 1313 -118
rect 1267 -1106 1273 -130
rect 1307 -1106 1313 -130
rect 1267 -1118 1313 -1106
rect 1525 -130 1571 -118
rect 1525 -1106 1531 -130
rect 1565 -1106 1571 -130
rect 1525 -1118 1571 -1106
rect 1783 -130 1829 -118
rect 1783 -1106 1789 -130
rect 1823 -1106 1829 -130
rect 1783 -1118 1829 -1106
rect 2041 -130 2087 -118
rect 2041 -1106 2047 -130
rect 2081 -1106 2087 -130
rect 2041 -1118 2087 -1106
rect 2299 -130 2345 -118
rect 2299 -1106 2305 -130
rect 2339 -1106 2345 -130
rect 2299 -1118 2345 -1106
rect 2557 -130 2603 -118
rect 2557 -1106 2563 -130
rect 2597 -1106 2603 -130
rect 2557 -1118 2603 -1106
rect 2815 -130 2861 -118
rect 2815 -1106 2821 -130
rect 2855 -1106 2861 -130
rect 2815 -1118 2861 -1106
rect 3073 -130 3119 -118
rect 3073 -1106 3079 -130
rect 3113 -1106 3119 -130
rect 3073 -1118 3119 -1106
rect 3331 -130 3377 -118
rect 3331 -1106 3337 -130
rect 3371 -1106 3377 -130
rect 3331 -1118 3377 -1106
rect 3589 -130 3635 -118
rect 3589 -1106 3595 -130
rect 3629 -1106 3635 -130
rect 3589 -1118 3635 -1106
rect -3579 -1165 -3387 -1159
rect -3579 -1199 -3567 -1165
rect -3399 -1199 -3387 -1165
rect -3579 -1205 -3387 -1199
rect -3321 -1165 -3129 -1159
rect -3321 -1199 -3309 -1165
rect -3141 -1199 -3129 -1165
rect -3321 -1205 -3129 -1199
rect -3063 -1165 -2871 -1159
rect -3063 -1199 -3051 -1165
rect -2883 -1199 -2871 -1165
rect -3063 -1205 -2871 -1199
rect -2805 -1165 -2613 -1159
rect -2805 -1199 -2793 -1165
rect -2625 -1199 -2613 -1165
rect -2805 -1205 -2613 -1199
rect -2547 -1165 -2355 -1159
rect -2547 -1199 -2535 -1165
rect -2367 -1199 -2355 -1165
rect -2547 -1205 -2355 -1199
rect -2289 -1165 -2097 -1159
rect -2289 -1199 -2277 -1165
rect -2109 -1199 -2097 -1165
rect -2289 -1205 -2097 -1199
rect -2031 -1165 -1839 -1159
rect -2031 -1199 -2019 -1165
rect -1851 -1199 -1839 -1165
rect -2031 -1205 -1839 -1199
rect -1773 -1165 -1581 -1159
rect -1773 -1199 -1761 -1165
rect -1593 -1199 -1581 -1165
rect -1773 -1205 -1581 -1199
rect -1515 -1165 -1323 -1159
rect -1515 -1199 -1503 -1165
rect -1335 -1199 -1323 -1165
rect -1515 -1205 -1323 -1199
rect -1257 -1165 -1065 -1159
rect -1257 -1199 -1245 -1165
rect -1077 -1199 -1065 -1165
rect -1257 -1205 -1065 -1199
rect -999 -1165 -807 -1159
rect -999 -1199 -987 -1165
rect -819 -1199 -807 -1165
rect -999 -1205 -807 -1199
rect -741 -1165 -549 -1159
rect -741 -1199 -729 -1165
rect -561 -1199 -549 -1165
rect -741 -1205 -549 -1199
rect -483 -1165 -291 -1159
rect -483 -1199 -471 -1165
rect -303 -1199 -291 -1165
rect -483 -1205 -291 -1199
rect -225 -1165 -33 -1159
rect -225 -1199 -213 -1165
rect -45 -1199 -33 -1165
rect -225 -1205 -33 -1199
rect 33 -1165 225 -1159
rect 33 -1199 45 -1165
rect 213 -1199 225 -1165
rect 33 -1205 225 -1199
rect 291 -1165 483 -1159
rect 291 -1199 303 -1165
rect 471 -1199 483 -1165
rect 291 -1205 483 -1199
rect 549 -1165 741 -1159
rect 549 -1199 561 -1165
rect 729 -1199 741 -1165
rect 549 -1205 741 -1199
rect 807 -1165 999 -1159
rect 807 -1199 819 -1165
rect 987 -1199 999 -1165
rect 807 -1205 999 -1199
rect 1065 -1165 1257 -1159
rect 1065 -1199 1077 -1165
rect 1245 -1199 1257 -1165
rect 1065 -1205 1257 -1199
rect 1323 -1165 1515 -1159
rect 1323 -1199 1335 -1165
rect 1503 -1199 1515 -1165
rect 1323 -1205 1515 -1199
rect 1581 -1165 1773 -1159
rect 1581 -1199 1593 -1165
rect 1761 -1199 1773 -1165
rect 1581 -1205 1773 -1199
rect 1839 -1165 2031 -1159
rect 1839 -1199 1851 -1165
rect 2019 -1199 2031 -1165
rect 1839 -1205 2031 -1199
rect 2097 -1165 2289 -1159
rect 2097 -1199 2109 -1165
rect 2277 -1199 2289 -1165
rect 2097 -1205 2289 -1199
rect 2355 -1165 2547 -1159
rect 2355 -1199 2367 -1165
rect 2535 -1199 2547 -1165
rect 2355 -1205 2547 -1199
rect 2613 -1165 2805 -1159
rect 2613 -1199 2625 -1165
rect 2793 -1199 2805 -1165
rect 2613 -1205 2805 -1199
rect 2871 -1165 3063 -1159
rect 2871 -1199 2883 -1165
rect 3051 -1199 3063 -1165
rect 2871 -1205 3063 -1199
rect 3129 -1165 3321 -1159
rect 3129 -1199 3141 -1165
rect 3309 -1199 3321 -1165
rect 3129 -1205 3321 -1199
rect 3387 -1165 3579 -1159
rect 3387 -1199 3399 -1165
rect 3567 -1199 3579 -1165
rect 3387 -1205 3579 -1199
rect -3579 -1273 -3387 -1267
rect -3579 -1307 -3567 -1273
rect -3399 -1307 -3387 -1273
rect -3579 -1313 -3387 -1307
rect -3321 -1273 -3129 -1267
rect -3321 -1307 -3309 -1273
rect -3141 -1307 -3129 -1273
rect -3321 -1313 -3129 -1307
rect -3063 -1273 -2871 -1267
rect -3063 -1307 -3051 -1273
rect -2883 -1307 -2871 -1273
rect -3063 -1313 -2871 -1307
rect -2805 -1273 -2613 -1267
rect -2805 -1307 -2793 -1273
rect -2625 -1307 -2613 -1273
rect -2805 -1313 -2613 -1307
rect -2547 -1273 -2355 -1267
rect -2547 -1307 -2535 -1273
rect -2367 -1307 -2355 -1273
rect -2547 -1313 -2355 -1307
rect -2289 -1273 -2097 -1267
rect -2289 -1307 -2277 -1273
rect -2109 -1307 -2097 -1273
rect -2289 -1313 -2097 -1307
rect -2031 -1273 -1839 -1267
rect -2031 -1307 -2019 -1273
rect -1851 -1307 -1839 -1273
rect -2031 -1313 -1839 -1307
rect -1773 -1273 -1581 -1267
rect -1773 -1307 -1761 -1273
rect -1593 -1307 -1581 -1273
rect -1773 -1313 -1581 -1307
rect -1515 -1273 -1323 -1267
rect -1515 -1307 -1503 -1273
rect -1335 -1307 -1323 -1273
rect -1515 -1313 -1323 -1307
rect -1257 -1273 -1065 -1267
rect -1257 -1307 -1245 -1273
rect -1077 -1307 -1065 -1273
rect -1257 -1313 -1065 -1307
rect -999 -1273 -807 -1267
rect -999 -1307 -987 -1273
rect -819 -1307 -807 -1273
rect -999 -1313 -807 -1307
rect -741 -1273 -549 -1267
rect -741 -1307 -729 -1273
rect -561 -1307 -549 -1273
rect -741 -1313 -549 -1307
rect -483 -1273 -291 -1267
rect -483 -1307 -471 -1273
rect -303 -1307 -291 -1273
rect -483 -1313 -291 -1307
rect -225 -1273 -33 -1267
rect -225 -1307 -213 -1273
rect -45 -1307 -33 -1273
rect -225 -1313 -33 -1307
rect 33 -1273 225 -1267
rect 33 -1307 45 -1273
rect 213 -1307 225 -1273
rect 33 -1313 225 -1307
rect 291 -1273 483 -1267
rect 291 -1307 303 -1273
rect 471 -1307 483 -1273
rect 291 -1313 483 -1307
rect 549 -1273 741 -1267
rect 549 -1307 561 -1273
rect 729 -1307 741 -1273
rect 549 -1313 741 -1307
rect 807 -1273 999 -1267
rect 807 -1307 819 -1273
rect 987 -1307 999 -1273
rect 807 -1313 999 -1307
rect 1065 -1273 1257 -1267
rect 1065 -1307 1077 -1273
rect 1245 -1307 1257 -1273
rect 1065 -1313 1257 -1307
rect 1323 -1273 1515 -1267
rect 1323 -1307 1335 -1273
rect 1503 -1307 1515 -1273
rect 1323 -1313 1515 -1307
rect 1581 -1273 1773 -1267
rect 1581 -1307 1593 -1273
rect 1761 -1307 1773 -1273
rect 1581 -1313 1773 -1307
rect 1839 -1273 2031 -1267
rect 1839 -1307 1851 -1273
rect 2019 -1307 2031 -1273
rect 1839 -1313 2031 -1307
rect 2097 -1273 2289 -1267
rect 2097 -1307 2109 -1273
rect 2277 -1307 2289 -1273
rect 2097 -1313 2289 -1307
rect 2355 -1273 2547 -1267
rect 2355 -1307 2367 -1273
rect 2535 -1307 2547 -1273
rect 2355 -1313 2547 -1307
rect 2613 -1273 2805 -1267
rect 2613 -1307 2625 -1273
rect 2793 -1307 2805 -1273
rect 2613 -1313 2805 -1307
rect 2871 -1273 3063 -1267
rect 2871 -1307 2883 -1273
rect 3051 -1307 3063 -1273
rect 2871 -1313 3063 -1307
rect 3129 -1273 3321 -1267
rect 3129 -1307 3141 -1273
rect 3309 -1307 3321 -1273
rect 3129 -1313 3321 -1307
rect 3387 -1273 3579 -1267
rect 3387 -1307 3399 -1273
rect 3567 -1307 3579 -1273
rect 3387 -1313 3579 -1307
rect -3635 -1366 -3589 -1354
rect -3635 -2342 -3629 -1366
rect -3595 -2342 -3589 -1366
rect -3635 -2354 -3589 -2342
rect -3377 -1366 -3331 -1354
rect -3377 -2342 -3371 -1366
rect -3337 -2342 -3331 -1366
rect -3377 -2354 -3331 -2342
rect -3119 -1366 -3073 -1354
rect -3119 -2342 -3113 -1366
rect -3079 -2342 -3073 -1366
rect -3119 -2354 -3073 -2342
rect -2861 -1366 -2815 -1354
rect -2861 -2342 -2855 -1366
rect -2821 -2342 -2815 -1366
rect -2861 -2354 -2815 -2342
rect -2603 -1366 -2557 -1354
rect -2603 -2342 -2597 -1366
rect -2563 -2342 -2557 -1366
rect -2603 -2354 -2557 -2342
rect -2345 -1366 -2299 -1354
rect -2345 -2342 -2339 -1366
rect -2305 -2342 -2299 -1366
rect -2345 -2354 -2299 -2342
rect -2087 -1366 -2041 -1354
rect -2087 -2342 -2081 -1366
rect -2047 -2342 -2041 -1366
rect -2087 -2354 -2041 -2342
rect -1829 -1366 -1783 -1354
rect -1829 -2342 -1823 -1366
rect -1789 -2342 -1783 -1366
rect -1829 -2354 -1783 -2342
rect -1571 -1366 -1525 -1354
rect -1571 -2342 -1565 -1366
rect -1531 -2342 -1525 -1366
rect -1571 -2354 -1525 -2342
rect -1313 -1366 -1267 -1354
rect -1313 -2342 -1307 -1366
rect -1273 -2342 -1267 -1366
rect -1313 -2354 -1267 -2342
rect -1055 -1366 -1009 -1354
rect -1055 -2342 -1049 -1366
rect -1015 -2342 -1009 -1366
rect -1055 -2354 -1009 -2342
rect -797 -1366 -751 -1354
rect -797 -2342 -791 -1366
rect -757 -2342 -751 -1366
rect -797 -2354 -751 -2342
rect -539 -1366 -493 -1354
rect -539 -2342 -533 -1366
rect -499 -2342 -493 -1366
rect -539 -2354 -493 -2342
rect -281 -1366 -235 -1354
rect -281 -2342 -275 -1366
rect -241 -2342 -235 -1366
rect -281 -2354 -235 -2342
rect -23 -1366 23 -1354
rect -23 -2342 -17 -1366
rect 17 -2342 23 -1366
rect -23 -2354 23 -2342
rect 235 -1366 281 -1354
rect 235 -2342 241 -1366
rect 275 -2342 281 -1366
rect 235 -2354 281 -2342
rect 493 -1366 539 -1354
rect 493 -2342 499 -1366
rect 533 -2342 539 -1366
rect 493 -2354 539 -2342
rect 751 -1366 797 -1354
rect 751 -2342 757 -1366
rect 791 -2342 797 -1366
rect 751 -2354 797 -2342
rect 1009 -1366 1055 -1354
rect 1009 -2342 1015 -1366
rect 1049 -2342 1055 -1366
rect 1009 -2354 1055 -2342
rect 1267 -1366 1313 -1354
rect 1267 -2342 1273 -1366
rect 1307 -2342 1313 -1366
rect 1267 -2354 1313 -2342
rect 1525 -1366 1571 -1354
rect 1525 -2342 1531 -1366
rect 1565 -2342 1571 -1366
rect 1525 -2354 1571 -2342
rect 1783 -1366 1829 -1354
rect 1783 -2342 1789 -1366
rect 1823 -2342 1829 -1366
rect 1783 -2354 1829 -2342
rect 2041 -1366 2087 -1354
rect 2041 -2342 2047 -1366
rect 2081 -2342 2087 -1366
rect 2041 -2354 2087 -2342
rect 2299 -1366 2345 -1354
rect 2299 -2342 2305 -1366
rect 2339 -2342 2345 -1366
rect 2299 -2354 2345 -2342
rect 2557 -1366 2603 -1354
rect 2557 -2342 2563 -1366
rect 2597 -2342 2603 -1366
rect 2557 -2354 2603 -2342
rect 2815 -1366 2861 -1354
rect 2815 -2342 2821 -1366
rect 2855 -2342 2861 -1366
rect 2815 -2354 2861 -2342
rect 3073 -1366 3119 -1354
rect 3073 -2342 3079 -1366
rect 3113 -2342 3119 -1366
rect 3073 -2354 3119 -2342
rect 3331 -1366 3377 -1354
rect 3331 -2342 3337 -1366
rect 3371 -2342 3377 -1366
rect 3331 -2354 3377 -2342
rect 3589 -1366 3635 -1354
rect 3589 -2342 3595 -1366
rect 3629 -2342 3635 -1366
rect 3589 -2354 3635 -2342
rect -3579 -2401 -3387 -2395
rect -3579 -2435 -3567 -2401
rect -3399 -2435 -3387 -2401
rect -3579 -2441 -3387 -2435
rect -3321 -2401 -3129 -2395
rect -3321 -2435 -3309 -2401
rect -3141 -2435 -3129 -2401
rect -3321 -2441 -3129 -2435
rect -3063 -2401 -2871 -2395
rect -3063 -2435 -3051 -2401
rect -2883 -2435 -2871 -2401
rect -3063 -2441 -2871 -2435
rect -2805 -2401 -2613 -2395
rect -2805 -2435 -2793 -2401
rect -2625 -2435 -2613 -2401
rect -2805 -2441 -2613 -2435
rect -2547 -2401 -2355 -2395
rect -2547 -2435 -2535 -2401
rect -2367 -2435 -2355 -2401
rect -2547 -2441 -2355 -2435
rect -2289 -2401 -2097 -2395
rect -2289 -2435 -2277 -2401
rect -2109 -2435 -2097 -2401
rect -2289 -2441 -2097 -2435
rect -2031 -2401 -1839 -2395
rect -2031 -2435 -2019 -2401
rect -1851 -2435 -1839 -2401
rect -2031 -2441 -1839 -2435
rect -1773 -2401 -1581 -2395
rect -1773 -2435 -1761 -2401
rect -1593 -2435 -1581 -2401
rect -1773 -2441 -1581 -2435
rect -1515 -2401 -1323 -2395
rect -1515 -2435 -1503 -2401
rect -1335 -2435 -1323 -2401
rect -1515 -2441 -1323 -2435
rect -1257 -2401 -1065 -2395
rect -1257 -2435 -1245 -2401
rect -1077 -2435 -1065 -2401
rect -1257 -2441 -1065 -2435
rect -999 -2401 -807 -2395
rect -999 -2435 -987 -2401
rect -819 -2435 -807 -2401
rect -999 -2441 -807 -2435
rect -741 -2401 -549 -2395
rect -741 -2435 -729 -2401
rect -561 -2435 -549 -2401
rect -741 -2441 -549 -2435
rect -483 -2401 -291 -2395
rect -483 -2435 -471 -2401
rect -303 -2435 -291 -2401
rect -483 -2441 -291 -2435
rect -225 -2401 -33 -2395
rect -225 -2435 -213 -2401
rect -45 -2435 -33 -2401
rect -225 -2441 -33 -2435
rect 33 -2401 225 -2395
rect 33 -2435 45 -2401
rect 213 -2435 225 -2401
rect 33 -2441 225 -2435
rect 291 -2401 483 -2395
rect 291 -2435 303 -2401
rect 471 -2435 483 -2401
rect 291 -2441 483 -2435
rect 549 -2401 741 -2395
rect 549 -2435 561 -2401
rect 729 -2435 741 -2401
rect 549 -2441 741 -2435
rect 807 -2401 999 -2395
rect 807 -2435 819 -2401
rect 987 -2435 999 -2401
rect 807 -2441 999 -2435
rect 1065 -2401 1257 -2395
rect 1065 -2435 1077 -2401
rect 1245 -2435 1257 -2401
rect 1065 -2441 1257 -2435
rect 1323 -2401 1515 -2395
rect 1323 -2435 1335 -2401
rect 1503 -2435 1515 -2401
rect 1323 -2441 1515 -2435
rect 1581 -2401 1773 -2395
rect 1581 -2435 1593 -2401
rect 1761 -2435 1773 -2401
rect 1581 -2441 1773 -2435
rect 1839 -2401 2031 -2395
rect 1839 -2435 1851 -2401
rect 2019 -2435 2031 -2401
rect 1839 -2441 2031 -2435
rect 2097 -2401 2289 -2395
rect 2097 -2435 2109 -2401
rect 2277 -2435 2289 -2401
rect 2097 -2441 2289 -2435
rect 2355 -2401 2547 -2395
rect 2355 -2435 2367 -2401
rect 2535 -2435 2547 -2401
rect 2355 -2441 2547 -2435
rect 2613 -2401 2805 -2395
rect 2613 -2435 2625 -2401
rect 2793 -2435 2805 -2401
rect 2613 -2441 2805 -2435
rect 2871 -2401 3063 -2395
rect 2871 -2435 2883 -2401
rect 3051 -2435 3063 -2401
rect 2871 -2441 3063 -2435
rect 3129 -2401 3321 -2395
rect 3129 -2435 3141 -2401
rect 3309 -2435 3321 -2401
rect 3129 -2441 3321 -2435
rect 3387 -2401 3579 -2395
rect 3387 -2435 3399 -2401
rect 3567 -2435 3579 -2401
rect 3387 -2441 3579 -2435
<< properties >>
string FIXED_BBOX -3746 -2556 3746 2556
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 1 m 4 nf 28 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
