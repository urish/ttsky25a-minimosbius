magic
tech sky130A
magscale 1 2
timestamp 1757105855
<< pwell >>
rect -2411 -1367 2411 1367
<< mvnmos >>
rect -2183 109 -2083 1109
rect -2025 109 -1925 1109
rect -1867 109 -1767 1109
rect -1709 109 -1609 1109
rect -1551 109 -1451 1109
rect -1393 109 -1293 1109
rect -1235 109 -1135 1109
rect -1077 109 -977 1109
rect -919 109 -819 1109
rect -761 109 -661 1109
rect -603 109 -503 1109
rect -445 109 -345 1109
rect -287 109 -187 1109
rect -129 109 -29 1109
rect 29 109 129 1109
rect 187 109 287 1109
rect 345 109 445 1109
rect 503 109 603 1109
rect 661 109 761 1109
rect 819 109 919 1109
rect 977 109 1077 1109
rect 1135 109 1235 1109
rect 1293 109 1393 1109
rect 1451 109 1551 1109
rect 1609 109 1709 1109
rect 1767 109 1867 1109
rect 1925 109 2025 1109
rect 2083 109 2183 1109
rect -2183 -1109 -2083 -109
rect -2025 -1109 -1925 -109
rect -1867 -1109 -1767 -109
rect -1709 -1109 -1609 -109
rect -1551 -1109 -1451 -109
rect -1393 -1109 -1293 -109
rect -1235 -1109 -1135 -109
rect -1077 -1109 -977 -109
rect -919 -1109 -819 -109
rect -761 -1109 -661 -109
rect -603 -1109 -503 -109
rect -445 -1109 -345 -109
rect -287 -1109 -187 -109
rect -129 -1109 -29 -109
rect 29 -1109 129 -109
rect 187 -1109 287 -109
rect 345 -1109 445 -109
rect 503 -1109 603 -109
rect 661 -1109 761 -109
rect 819 -1109 919 -109
rect 977 -1109 1077 -109
rect 1135 -1109 1235 -109
rect 1293 -1109 1393 -109
rect 1451 -1109 1551 -109
rect 1609 -1109 1709 -109
rect 1767 -1109 1867 -109
rect 1925 -1109 2025 -109
rect 2083 -1109 2183 -109
<< mvndiff >>
rect -2241 1097 -2183 1109
rect -2241 121 -2229 1097
rect -2195 121 -2183 1097
rect -2241 109 -2183 121
rect -2083 1097 -2025 1109
rect -2083 121 -2071 1097
rect -2037 121 -2025 1097
rect -2083 109 -2025 121
rect -1925 1097 -1867 1109
rect -1925 121 -1913 1097
rect -1879 121 -1867 1097
rect -1925 109 -1867 121
rect -1767 1097 -1709 1109
rect -1767 121 -1755 1097
rect -1721 121 -1709 1097
rect -1767 109 -1709 121
rect -1609 1097 -1551 1109
rect -1609 121 -1597 1097
rect -1563 121 -1551 1097
rect -1609 109 -1551 121
rect -1451 1097 -1393 1109
rect -1451 121 -1439 1097
rect -1405 121 -1393 1097
rect -1451 109 -1393 121
rect -1293 1097 -1235 1109
rect -1293 121 -1281 1097
rect -1247 121 -1235 1097
rect -1293 109 -1235 121
rect -1135 1097 -1077 1109
rect -1135 121 -1123 1097
rect -1089 121 -1077 1097
rect -1135 109 -1077 121
rect -977 1097 -919 1109
rect -977 121 -965 1097
rect -931 121 -919 1097
rect -977 109 -919 121
rect -819 1097 -761 1109
rect -819 121 -807 1097
rect -773 121 -761 1097
rect -819 109 -761 121
rect -661 1097 -603 1109
rect -661 121 -649 1097
rect -615 121 -603 1097
rect -661 109 -603 121
rect -503 1097 -445 1109
rect -503 121 -491 1097
rect -457 121 -445 1097
rect -503 109 -445 121
rect -345 1097 -287 1109
rect -345 121 -333 1097
rect -299 121 -287 1097
rect -345 109 -287 121
rect -187 1097 -129 1109
rect -187 121 -175 1097
rect -141 121 -129 1097
rect -187 109 -129 121
rect -29 1097 29 1109
rect -29 121 -17 1097
rect 17 121 29 1097
rect -29 109 29 121
rect 129 1097 187 1109
rect 129 121 141 1097
rect 175 121 187 1097
rect 129 109 187 121
rect 287 1097 345 1109
rect 287 121 299 1097
rect 333 121 345 1097
rect 287 109 345 121
rect 445 1097 503 1109
rect 445 121 457 1097
rect 491 121 503 1097
rect 445 109 503 121
rect 603 1097 661 1109
rect 603 121 615 1097
rect 649 121 661 1097
rect 603 109 661 121
rect 761 1097 819 1109
rect 761 121 773 1097
rect 807 121 819 1097
rect 761 109 819 121
rect 919 1097 977 1109
rect 919 121 931 1097
rect 965 121 977 1097
rect 919 109 977 121
rect 1077 1097 1135 1109
rect 1077 121 1089 1097
rect 1123 121 1135 1097
rect 1077 109 1135 121
rect 1235 1097 1293 1109
rect 1235 121 1247 1097
rect 1281 121 1293 1097
rect 1235 109 1293 121
rect 1393 1097 1451 1109
rect 1393 121 1405 1097
rect 1439 121 1451 1097
rect 1393 109 1451 121
rect 1551 1097 1609 1109
rect 1551 121 1563 1097
rect 1597 121 1609 1097
rect 1551 109 1609 121
rect 1709 1097 1767 1109
rect 1709 121 1721 1097
rect 1755 121 1767 1097
rect 1709 109 1767 121
rect 1867 1097 1925 1109
rect 1867 121 1879 1097
rect 1913 121 1925 1097
rect 1867 109 1925 121
rect 2025 1097 2083 1109
rect 2025 121 2037 1097
rect 2071 121 2083 1097
rect 2025 109 2083 121
rect 2183 1097 2241 1109
rect 2183 121 2195 1097
rect 2229 121 2241 1097
rect 2183 109 2241 121
rect -2241 -121 -2183 -109
rect -2241 -1097 -2229 -121
rect -2195 -1097 -2183 -121
rect -2241 -1109 -2183 -1097
rect -2083 -121 -2025 -109
rect -2083 -1097 -2071 -121
rect -2037 -1097 -2025 -121
rect -2083 -1109 -2025 -1097
rect -1925 -121 -1867 -109
rect -1925 -1097 -1913 -121
rect -1879 -1097 -1867 -121
rect -1925 -1109 -1867 -1097
rect -1767 -121 -1709 -109
rect -1767 -1097 -1755 -121
rect -1721 -1097 -1709 -121
rect -1767 -1109 -1709 -1097
rect -1609 -121 -1551 -109
rect -1609 -1097 -1597 -121
rect -1563 -1097 -1551 -121
rect -1609 -1109 -1551 -1097
rect -1451 -121 -1393 -109
rect -1451 -1097 -1439 -121
rect -1405 -1097 -1393 -121
rect -1451 -1109 -1393 -1097
rect -1293 -121 -1235 -109
rect -1293 -1097 -1281 -121
rect -1247 -1097 -1235 -121
rect -1293 -1109 -1235 -1097
rect -1135 -121 -1077 -109
rect -1135 -1097 -1123 -121
rect -1089 -1097 -1077 -121
rect -1135 -1109 -1077 -1097
rect -977 -121 -919 -109
rect -977 -1097 -965 -121
rect -931 -1097 -919 -121
rect -977 -1109 -919 -1097
rect -819 -121 -761 -109
rect -819 -1097 -807 -121
rect -773 -1097 -761 -121
rect -819 -1109 -761 -1097
rect -661 -121 -603 -109
rect -661 -1097 -649 -121
rect -615 -1097 -603 -121
rect -661 -1109 -603 -1097
rect -503 -121 -445 -109
rect -503 -1097 -491 -121
rect -457 -1097 -445 -121
rect -503 -1109 -445 -1097
rect -345 -121 -287 -109
rect -345 -1097 -333 -121
rect -299 -1097 -287 -121
rect -345 -1109 -287 -1097
rect -187 -121 -129 -109
rect -187 -1097 -175 -121
rect -141 -1097 -129 -121
rect -187 -1109 -129 -1097
rect -29 -121 29 -109
rect -29 -1097 -17 -121
rect 17 -1097 29 -121
rect -29 -1109 29 -1097
rect 129 -121 187 -109
rect 129 -1097 141 -121
rect 175 -1097 187 -121
rect 129 -1109 187 -1097
rect 287 -121 345 -109
rect 287 -1097 299 -121
rect 333 -1097 345 -121
rect 287 -1109 345 -1097
rect 445 -121 503 -109
rect 445 -1097 457 -121
rect 491 -1097 503 -121
rect 445 -1109 503 -1097
rect 603 -121 661 -109
rect 603 -1097 615 -121
rect 649 -1097 661 -121
rect 603 -1109 661 -1097
rect 761 -121 819 -109
rect 761 -1097 773 -121
rect 807 -1097 819 -121
rect 761 -1109 819 -1097
rect 919 -121 977 -109
rect 919 -1097 931 -121
rect 965 -1097 977 -121
rect 919 -1109 977 -1097
rect 1077 -121 1135 -109
rect 1077 -1097 1089 -121
rect 1123 -1097 1135 -121
rect 1077 -1109 1135 -1097
rect 1235 -121 1293 -109
rect 1235 -1097 1247 -121
rect 1281 -1097 1293 -121
rect 1235 -1109 1293 -1097
rect 1393 -121 1451 -109
rect 1393 -1097 1405 -121
rect 1439 -1097 1451 -121
rect 1393 -1109 1451 -1097
rect 1551 -121 1609 -109
rect 1551 -1097 1563 -121
rect 1597 -1097 1609 -121
rect 1551 -1109 1609 -1097
rect 1709 -121 1767 -109
rect 1709 -1097 1721 -121
rect 1755 -1097 1767 -121
rect 1709 -1109 1767 -1097
rect 1867 -121 1925 -109
rect 1867 -1097 1879 -121
rect 1913 -1097 1925 -121
rect 1867 -1109 1925 -1097
rect 2025 -121 2083 -109
rect 2025 -1097 2037 -121
rect 2071 -1097 2083 -121
rect 2025 -1109 2083 -1097
rect 2183 -121 2241 -109
rect 2183 -1097 2195 -121
rect 2229 -1097 2241 -121
rect 2183 -1109 2241 -1097
<< mvndiffc >>
rect -2229 121 -2195 1097
rect -2071 121 -2037 1097
rect -1913 121 -1879 1097
rect -1755 121 -1721 1097
rect -1597 121 -1563 1097
rect -1439 121 -1405 1097
rect -1281 121 -1247 1097
rect -1123 121 -1089 1097
rect -965 121 -931 1097
rect -807 121 -773 1097
rect -649 121 -615 1097
rect -491 121 -457 1097
rect -333 121 -299 1097
rect -175 121 -141 1097
rect -17 121 17 1097
rect 141 121 175 1097
rect 299 121 333 1097
rect 457 121 491 1097
rect 615 121 649 1097
rect 773 121 807 1097
rect 931 121 965 1097
rect 1089 121 1123 1097
rect 1247 121 1281 1097
rect 1405 121 1439 1097
rect 1563 121 1597 1097
rect 1721 121 1755 1097
rect 1879 121 1913 1097
rect 2037 121 2071 1097
rect 2195 121 2229 1097
rect -2229 -1097 -2195 -121
rect -2071 -1097 -2037 -121
rect -1913 -1097 -1879 -121
rect -1755 -1097 -1721 -121
rect -1597 -1097 -1563 -121
rect -1439 -1097 -1405 -121
rect -1281 -1097 -1247 -121
rect -1123 -1097 -1089 -121
rect -965 -1097 -931 -121
rect -807 -1097 -773 -121
rect -649 -1097 -615 -121
rect -491 -1097 -457 -121
rect -333 -1097 -299 -121
rect -175 -1097 -141 -121
rect -17 -1097 17 -121
rect 141 -1097 175 -121
rect 299 -1097 333 -121
rect 457 -1097 491 -121
rect 615 -1097 649 -121
rect 773 -1097 807 -121
rect 931 -1097 965 -121
rect 1089 -1097 1123 -121
rect 1247 -1097 1281 -121
rect 1405 -1097 1439 -121
rect 1563 -1097 1597 -121
rect 1721 -1097 1755 -121
rect 1879 -1097 1913 -121
rect 2037 -1097 2071 -121
rect 2195 -1097 2229 -121
<< mvpsubdiff >>
rect -2375 1319 2375 1331
rect -2375 1285 -2267 1319
rect 2267 1285 2375 1319
rect -2375 1273 2375 1285
rect -2375 1223 -2317 1273
rect -2375 -1223 -2363 1223
rect -2329 -1223 -2317 1223
rect 2317 1223 2375 1273
rect -2375 -1273 -2317 -1223
rect 2317 -1223 2329 1223
rect 2363 -1223 2375 1223
rect 2317 -1273 2375 -1223
rect -2375 -1285 2375 -1273
rect -2375 -1319 -2267 -1285
rect 2267 -1319 2375 -1285
rect -2375 -1331 2375 -1319
<< mvpsubdiffcont >>
rect -2267 1285 2267 1319
rect -2363 -1223 -2329 1223
rect 2329 -1223 2363 1223
rect -2267 -1319 2267 -1285
<< poly >>
rect -2183 1181 -2083 1197
rect -2183 1147 -2167 1181
rect -2099 1147 -2083 1181
rect -2183 1109 -2083 1147
rect -2025 1181 -1925 1197
rect -2025 1147 -2009 1181
rect -1941 1147 -1925 1181
rect -2025 1109 -1925 1147
rect -1867 1181 -1767 1197
rect -1867 1147 -1851 1181
rect -1783 1147 -1767 1181
rect -1867 1109 -1767 1147
rect -1709 1181 -1609 1197
rect -1709 1147 -1693 1181
rect -1625 1147 -1609 1181
rect -1709 1109 -1609 1147
rect -1551 1181 -1451 1197
rect -1551 1147 -1535 1181
rect -1467 1147 -1451 1181
rect -1551 1109 -1451 1147
rect -1393 1181 -1293 1197
rect -1393 1147 -1377 1181
rect -1309 1147 -1293 1181
rect -1393 1109 -1293 1147
rect -1235 1181 -1135 1197
rect -1235 1147 -1219 1181
rect -1151 1147 -1135 1181
rect -1235 1109 -1135 1147
rect -1077 1181 -977 1197
rect -1077 1147 -1061 1181
rect -993 1147 -977 1181
rect -1077 1109 -977 1147
rect -919 1181 -819 1197
rect -919 1147 -903 1181
rect -835 1147 -819 1181
rect -919 1109 -819 1147
rect -761 1181 -661 1197
rect -761 1147 -745 1181
rect -677 1147 -661 1181
rect -761 1109 -661 1147
rect -603 1181 -503 1197
rect -603 1147 -587 1181
rect -519 1147 -503 1181
rect -603 1109 -503 1147
rect -445 1181 -345 1197
rect -445 1147 -429 1181
rect -361 1147 -345 1181
rect -445 1109 -345 1147
rect -287 1181 -187 1197
rect -287 1147 -271 1181
rect -203 1147 -187 1181
rect -287 1109 -187 1147
rect -129 1181 -29 1197
rect -129 1147 -113 1181
rect -45 1147 -29 1181
rect -129 1109 -29 1147
rect 29 1181 129 1197
rect 29 1147 45 1181
rect 113 1147 129 1181
rect 29 1109 129 1147
rect 187 1181 287 1197
rect 187 1147 203 1181
rect 271 1147 287 1181
rect 187 1109 287 1147
rect 345 1181 445 1197
rect 345 1147 361 1181
rect 429 1147 445 1181
rect 345 1109 445 1147
rect 503 1181 603 1197
rect 503 1147 519 1181
rect 587 1147 603 1181
rect 503 1109 603 1147
rect 661 1181 761 1197
rect 661 1147 677 1181
rect 745 1147 761 1181
rect 661 1109 761 1147
rect 819 1181 919 1197
rect 819 1147 835 1181
rect 903 1147 919 1181
rect 819 1109 919 1147
rect 977 1181 1077 1197
rect 977 1147 993 1181
rect 1061 1147 1077 1181
rect 977 1109 1077 1147
rect 1135 1181 1235 1197
rect 1135 1147 1151 1181
rect 1219 1147 1235 1181
rect 1135 1109 1235 1147
rect 1293 1181 1393 1197
rect 1293 1147 1309 1181
rect 1377 1147 1393 1181
rect 1293 1109 1393 1147
rect 1451 1181 1551 1197
rect 1451 1147 1467 1181
rect 1535 1147 1551 1181
rect 1451 1109 1551 1147
rect 1609 1181 1709 1197
rect 1609 1147 1625 1181
rect 1693 1147 1709 1181
rect 1609 1109 1709 1147
rect 1767 1181 1867 1197
rect 1767 1147 1783 1181
rect 1851 1147 1867 1181
rect 1767 1109 1867 1147
rect 1925 1181 2025 1197
rect 1925 1147 1941 1181
rect 2009 1147 2025 1181
rect 1925 1109 2025 1147
rect 2083 1181 2183 1197
rect 2083 1147 2099 1181
rect 2167 1147 2183 1181
rect 2083 1109 2183 1147
rect -2183 71 -2083 109
rect -2183 37 -2167 71
rect -2099 37 -2083 71
rect -2183 21 -2083 37
rect -2025 71 -1925 109
rect -2025 37 -2009 71
rect -1941 37 -1925 71
rect -2025 21 -1925 37
rect -1867 71 -1767 109
rect -1867 37 -1851 71
rect -1783 37 -1767 71
rect -1867 21 -1767 37
rect -1709 71 -1609 109
rect -1709 37 -1693 71
rect -1625 37 -1609 71
rect -1709 21 -1609 37
rect -1551 71 -1451 109
rect -1551 37 -1535 71
rect -1467 37 -1451 71
rect -1551 21 -1451 37
rect -1393 71 -1293 109
rect -1393 37 -1377 71
rect -1309 37 -1293 71
rect -1393 21 -1293 37
rect -1235 71 -1135 109
rect -1235 37 -1219 71
rect -1151 37 -1135 71
rect -1235 21 -1135 37
rect -1077 71 -977 109
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -1077 21 -977 37
rect -919 71 -819 109
rect -919 37 -903 71
rect -835 37 -819 71
rect -919 21 -819 37
rect -761 71 -661 109
rect -761 37 -745 71
rect -677 37 -661 71
rect -761 21 -661 37
rect -603 71 -503 109
rect -603 37 -587 71
rect -519 37 -503 71
rect -603 21 -503 37
rect -445 71 -345 109
rect -445 37 -429 71
rect -361 37 -345 71
rect -445 21 -345 37
rect -287 71 -187 109
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 109
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 109
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 109
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect 345 71 445 109
rect 345 37 361 71
rect 429 37 445 71
rect 345 21 445 37
rect 503 71 603 109
rect 503 37 519 71
rect 587 37 603 71
rect 503 21 603 37
rect 661 71 761 109
rect 661 37 677 71
rect 745 37 761 71
rect 661 21 761 37
rect 819 71 919 109
rect 819 37 835 71
rect 903 37 919 71
rect 819 21 919 37
rect 977 71 1077 109
rect 977 37 993 71
rect 1061 37 1077 71
rect 977 21 1077 37
rect 1135 71 1235 109
rect 1135 37 1151 71
rect 1219 37 1235 71
rect 1135 21 1235 37
rect 1293 71 1393 109
rect 1293 37 1309 71
rect 1377 37 1393 71
rect 1293 21 1393 37
rect 1451 71 1551 109
rect 1451 37 1467 71
rect 1535 37 1551 71
rect 1451 21 1551 37
rect 1609 71 1709 109
rect 1609 37 1625 71
rect 1693 37 1709 71
rect 1609 21 1709 37
rect 1767 71 1867 109
rect 1767 37 1783 71
rect 1851 37 1867 71
rect 1767 21 1867 37
rect 1925 71 2025 109
rect 1925 37 1941 71
rect 2009 37 2025 71
rect 1925 21 2025 37
rect 2083 71 2183 109
rect 2083 37 2099 71
rect 2167 37 2183 71
rect 2083 21 2183 37
rect -2183 -37 -2083 -21
rect -2183 -71 -2167 -37
rect -2099 -71 -2083 -37
rect -2183 -109 -2083 -71
rect -2025 -37 -1925 -21
rect -2025 -71 -2009 -37
rect -1941 -71 -1925 -37
rect -2025 -109 -1925 -71
rect -1867 -37 -1767 -21
rect -1867 -71 -1851 -37
rect -1783 -71 -1767 -37
rect -1867 -109 -1767 -71
rect -1709 -37 -1609 -21
rect -1709 -71 -1693 -37
rect -1625 -71 -1609 -37
rect -1709 -109 -1609 -71
rect -1551 -37 -1451 -21
rect -1551 -71 -1535 -37
rect -1467 -71 -1451 -37
rect -1551 -109 -1451 -71
rect -1393 -37 -1293 -21
rect -1393 -71 -1377 -37
rect -1309 -71 -1293 -37
rect -1393 -109 -1293 -71
rect -1235 -37 -1135 -21
rect -1235 -71 -1219 -37
rect -1151 -71 -1135 -37
rect -1235 -109 -1135 -71
rect -1077 -37 -977 -21
rect -1077 -71 -1061 -37
rect -993 -71 -977 -37
rect -1077 -109 -977 -71
rect -919 -37 -819 -21
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -919 -109 -819 -71
rect -761 -37 -661 -21
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -761 -109 -661 -71
rect -603 -37 -503 -21
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -603 -109 -503 -71
rect -445 -37 -345 -21
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -445 -109 -345 -71
rect -287 -37 -187 -21
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -287 -109 -187 -71
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -109 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -109 129 -71
rect 187 -37 287 -21
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 187 -109 287 -71
rect 345 -37 445 -21
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 345 -109 445 -71
rect 503 -37 603 -21
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 503 -109 603 -71
rect 661 -37 761 -21
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 661 -109 761 -71
rect 819 -37 919 -21
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 819 -109 919 -71
rect 977 -37 1077 -21
rect 977 -71 993 -37
rect 1061 -71 1077 -37
rect 977 -109 1077 -71
rect 1135 -37 1235 -21
rect 1135 -71 1151 -37
rect 1219 -71 1235 -37
rect 1135 -109 1235 -71
rect 1293 -37 1393 -21
rect 1293 -71 1309 -37
rect 1377 -71 1393 -37
rect 1293 -109 1393 -71
rect 1451 -37 1551 -21
rect 1451 -71 1467 -37
rect 1535 -71 1551 -37
rect 1451 -109 1551 -71
rect 1609 -37 1709 -21
rect 1609 -71 1625 -37
rect 1693 -71 1709 -37
rect 1609 -109 1709 -71
rect 1767 -37 1867 -21
rect 1767 -71 1783 -37
rect 1851 -71 1867 -37
rect 1767 -109 1867 -71
rect 1925 -37 2025 -21
rect 1925 -71 1941 -37
rect 2009 -71 2025 -37
rect 1925 -109 2025 -71
rect 2083 -37 2183 -21
rect 2083 -71 2099 -37
rect 2167 -71 2183 -37
rect 2083 -109 2183 -71
rect -2183 -1147 -2083 -1109
rect -2183 -1181 -2167 -1147
rect -2099 -1181 -2083 -1147
rect -2183 -1197 -2083 -1181
rect -2025 -1147 -1925 -1109
rect -2025 -1181 -2009 -1147
rect -1941 -1181 -1925 -1147
rect -2025 -1197 -1925 -1181
rect -1867 -1147 -1767 -1109
rect -1867 -1181 -1851 -1147
rect -1783 -1181 -1767 -1147
rect -1867 -1197 -1767 -1181
rect -1709 -1147 -1609 -1109
rect -1709 -1181 -1693 -1147
rect -1625 -1181 -1609 -1147
rect -1709 -1197 -1609 -1181
rect -1551 -1147 -1451 -1109
rect -1551 -1181 -1535 -1147
rect -1467 -1181 -1451 -1147
rect -1551 -1197 -1451 -1181
rect -1393 -1147 -1293 -1109
rect -1393 -1181 -1377 -1147
rect -1309 -1181 -1293 -1147
rect -1393 -1197 -1293 -1181
rect -1235 -1147 -1135 -1109
rect -1235 -1181 -1219 -1147
rect -1151 -1181 -1135 -1147
rect -1235 -1197 -1135 -1181
rect -1077 -1147 -977 -1109
rect -1077 -1181 -1061 -1147
rect -993 -1181 -977 -1147
rect -1077 -1197 -977 -1181
rect -919 -1147 -819 -1109
rect -919 -1181 -903 -1147
rect -835 -1181 -819 -1147
rect -919 -1197 -819 -1181
rect -761 -1147 -661 -1109
rect -761 -1181 -745 -1147
rect -677 -1181 -661 -1147
rect -761 -1197 -661 -1181
rect -603 -1147 -503 -1109
rect -603 -1181 -587 -1147
rect -519 -1181 -503 -1147
rect -603 -1197 -503 -1181
rect -445 -1147 -345 -1109
rect -445 -1181 -429 -1147
rect -361 -1181 -345 -1147
rect -445 -1197 -345 -1181
rect -287 -1147 -187 -1109
rect -287 -1181 -271 -1147
rect -203 -1181 -187 -1147
rect -287 -1197 -187 -1181
rect -129 -1147 -29 -1109
rect -129 -1181 -113 -1147
rect -45 -1181 -29 -1147
rect -129 -1197 -29 -1181
rect 29 -1147 129 -1109
rect 29 -1181 45 -1147
rect 113 -1181 129 -1147
rect 29 -1197 129 -1181
rect 187 -1147 287 -1109
rect 187 -1181 203 -1147
rect 271 -1181 287 -1147
rect 187 -1197 287 -1181
rect 345 -1147 445 -1109
rect 345 -1181 361 -1147
rect 429 -1181 445 -1147
rect 345 -1197 445 -1181
rect 503 -1147 603 -1109
rect 503 -1181 519 -1147
rect 587 -1181 603 -1147
rect 503 -1197 603 -1181
rect 661 -1147 761 -1109
rect 661 -1181 677 -1147
rect 745 -1181 761 -1147
rect 661 -1197 761 -1181
rect 819 -1147 919 -1109
rect 819 -1181 835 -1147
rect 903 -1181 919 -1147
rect 819 -1197 919 -1181
rect 977 -1147 1077 -1109
rect 977 -1181 993 -1147
rect 1061 -1181 1077 -1147
rect 977 -1197 1077 -1181
rect 1135 -1147 1235 -1109
rect 1135 -1181 1151 -1147
rect 1219 -1181 1235 -1147
rect 1135 -1197 1235 -1181
rect 1293 -1147 1393 -1109
rect 1293 -1181 1309 -1147
rect 1377 -1181 1393 -1147
rect 1293 -1197 1393 -1181
rect 1451 -1147 1551 -1109
rect 1451 -1181 1467 -1147
rect 1535 -1181 1551 -1147
rect 1451 -1197 1551 -1181
rect 1609 -1147 1709 -1109
rect 1609 -1181 1625 -1147
rect 1693 -1181 1709 -1147
rect 1609 -1197 1709 -1181
rect 1767 -1147 1867 -1109
rect 1767 -1181 1783 -1147
rect 1851 -1181 1867 -1147
rect 1767 -1197 1867 -1181
rect 1925 -1147 2025 -1109
rect 1925 -1181 1941 -1147
rect 2009 -1181 2025 -1147
rect 1925 -1197 2025 -1181
rect 2083 -1147 2183 -1109
rect 2083 -1181 2099 -1147
rect 2167 -1181 2183 -1147
rect 2083 -1197 2183 -1181
<< polycont >>
rect -2167 1147 -2099 1181
rect -2009 1147 -1941 1181
rect -1851 1147 -1783 1181
rect -1693 1147 -1625 1181
rect -1535 1147 -1467 1181
rect -1377 1147 -1309 1181
rect -1219 1147 -1151 1181
rect -1061 1147 -993 1181
rect -903 1147 -835 1181
rect -745 1147 -677 1181
rect -587 1147 -519 1181
rect -429 1147 -361 1181
rect -271 1147 -203 1181
rect -113 1147 -45 1181
rect 45 1147 113 1181
rect 203 1147 271 1181
rect 361 1147 429 1181
rect 519 1147 587 1181
rect 677 1147 745 1181
rect 835 1147 903 1181
rect 993 1147 1061 1181
rect 1151 1147 1219 1181
rect 1309 1147 1377 1181
rect 1467 1147 1535 1181
rect 1625 1147 1693 1181
rect 1783 1147 1851 1181
rect 1941 1147 2009 1181
rect 2099 1147 2167 1181
rect -2167 37 -2099 71
rect -2009 37 -1941 71
rect -1851 37 -1783 71
rect -1693 37 -1625 71
rect -1535 37 -1467 71
rect -1377 37 -1309 71
rect -1219 37 -1151 71
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect 1151 37 1219 71
rect 1309 37 1377 71
rect 1467 37 1535 71
rect 1625 37 1693 71
rect 1783 37 1851 71
rect 1941 37 2009 71
rect 2099 37 2167 71
rect -2167 -71 -2099 -37
rect -2009 -71 -1941 -37
rect -1851 -71 -1783 -37
rect -1693 -71 -1625 -37
rect -1535 -71 -1467 -37
rect -1377 -71 -1309 -37
rect -1219 -71 -1151 -37
rect -1061 -71 -993 -37
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect 993 -71 1061 -37
rect 1151 -71 1219 -37
rect 1309 -71 1377 -37
rect 1467 -71 1535 -37
rect 1625 -71 1693 -37
rect 1783 -71 1851 -37
rect 1941 -71 2009 -37
rect 2099 -71 2167 -37
rect -2167 -1181 -2099 -1147
rect -2009 -1181 -1941 -1147
rect -1851 -1181 -1783 -1147
rect -1693 -1181 -1625 -1147
rect -1535 -1181 -1467 -1147
rect -1377 -1181 -1309 -1147
rect -1219 -1181 -1151 -1147
rect -1061 -1181 -993 -1147
rect -903 -1181 -835 -1147
rect -745 -1181 -677 -1147
rect -587 -1181 -519 -1147
rect -429 -1181 -361 -1147
rect -271 -1181 -203 -1147
rect -113 -1181 -45 -1147
rect 45 -1181 113 -1147
rect 203 -1181 271 -1147
rect 361 -1181 429 -1147
rect 519 -1181 587 -1147
rect 677 -1181 745 -1147
rect 835 -1181 903 -1147
rect 993 -1181 1061 -1147
rect 1151 -1181 1219 -1147
rect 1309 -1181 1377 -1147
rect 1467 -1181 1535 -1147
rect 1625 -1181 1693 -1147
rect 1783 -1181 1851 -1147
rect 1941 -1181 2009 -1147
rect 2099 -1181 2167 -1147
<< locali >>
rect -2363 1285 -2267 1319
rect 2267 1285 2363 1319
rect -2363 1223 -2329 1285
rect 2329 1223 2363 1285
rect -2183 1147 -2167 1181
rect -2099 1147 -2083 1181
rect -2025 1147 -2009 1181
rect -1941 1147 -1925 1181
rect -1867 1147 -1851 1181
rect -1783 1147 -1767 1181
rect -1709 1147 -1693 1181
rect -1625 1147 -1609 1181
rect -1551 1147 -1535 1181
rect -1467 1147 -1451 1181
rect -1393 1147 -1377 1181
rect -1309 1147 -1293 1181
rect -1235 1147 -1219 1181
rect -1151 1147 -1135 1181
rect -1077 1147 -1061 1181
rect -993 1147 -977 1181
rect -919 1147 -903 1181
rect -835 1147 -819 1181
rect -761 1147 -745 1181
rect -677 1147 -661 1181
rect -603 1147 -587 1181
rect -519 1147 -503 1181
rect -445 1147 -429 1181
rect -361 1147 -345 1181
rect -287 1147 -271 1181
rect -203 1147 -187 1181
rect -129 1147 -113 1181
rect -45 1147 -29 1181
rect 29 1147 45 1181
rect 113 1147 129 1181
rect 187 1147 203 1181
rect 271 1147 287 1181
rect 345 1147 361 1181
rect 429 1147 445 1181
rect 503 1147 519 1181
rect 587 1147 603 1181
rect 661 1147 677 1181
rect 745 1147 761 1181
rect 819 1147 835 1181
rect 903 1147 919 1181
rect 977 1147 993 1181
rect 1061 1147 1077 1181
rect 1135 1147 1151 1181
rect 1219 1147 1235 1181
rect 1293 1147 1309 1181
rect 1377 1147 1393 1181
rect 1451 1147 1467 1181
rect 1535 1147 1551 1181
rect 1609 1147 1625 1181
rect 1693 1147 1709 1181
rect 1767 1147 1783 1181
rect 1851 1147 1867 1181
rect 1925 1147 1941 1181
rect 2009 1147 2025 1181
rect 2083 1147 2099 1181
rect 2167 1147 2183 1181
rect -2229 1097 -2195 1113
rect -2229 105 -2195 121
rect -2071 1097 -2037 1113
rect -2071 105 -2037 121
rect -1913 1097 -1879 1113
rect -1913 105 -1879 121
rect -1755 1097 -1721 1113
rect -1755 105 -1721 121
rect -1597 1097 -1563 1113
rect -1597 105 -1563 121
rect -1439 1097 -1405 1113
rect -1439 105 -1405 121
rect -1281 1097 -1247 1113
rect -1281 105 -1247 121
rect -1123 1097 -1089 1113
rect -1123 105 -1089 121
rect -965 1097 -931 1113
rect -965 105 -931 121
rect -807 1097 -773 1113
rect -807 105 -773 121
rect -649 1097 -615 1113
rect -649 105 -615 121
rect -491 1097 -457 1113
rect -491 105 -457 121
rect -333 1097 -299 1113
rect -333 105 -299 121
rect -175 1097 -141 1113
rect -175 105 -141 121
rect -17 1097 17 1113
rect -17 105 17 121
rect 141 1097 175 1113
rect 141 105 175 121
rect 299 1097 333 1113
rect 299 105 333 121
rect 457 1097 491 1113
rect 457 105 491 121
rect 615 1097 649 1113
rect 615 105 649 121
rect 773 1097 807 1113
rect 773 105 807 121
rect 931 1097 965 1113
rect 931 105 965 121
rect 1089 1097 1123 1113
rect 1089 105 1123 121
rect 1247 1097 1281 1113
rect 1247 105 1281 121
rect 1405 1097 1439 1113
rect 1405 105 1439 121
rect 1563 1097 1597 1113
rect 1563 105 1597 121
rect 1721 1097 1755 1113
rect 1721 105 1755 121
rect 1879 1097 1913 1113
rect 1879 105 1913 121
rect 2037 1097 2071 1113
rect 2037 105 2071 121
rect 2195 1097 2229 1113
rect 2195 105 2229 121
rect -2183 37 -2167 71
rect -2099 37 -2083 71
rect -2025 37 -2009 71
rect -1941 37 -1925 71
rect -1867 37 -1851 71
rect -1783 37 -1767 71
rect -1709 37 -1693 71
rect -1625 37 -1609 71
rect -1551 37 -1535 71
rect -1467 37 -1451 71
rect -1393 37 -1377 71
rect -1309 37 -1293 71
rect -1235 37 -1219 71
rect -1151 37 -1135 71
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -919 37 -903 71
rect -835 37 -819 71
rect -761 37 -745 71
rect -677 37 -661 71
rect -603 37 -587 71
rect -519 37 -503 71
rect -445 37 -429 71
rect -361 37 -345 71
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect 345 37 361 71
rect 429 37 445 71
rect 503 37 519 71
rect 587 37 603 71
rect 661 37 677 71
rect 745 37 761 71
rect 819 37 835 71
rect 903 37 919 71
rect 977 37 993 71
rect 1061 37 1077 71
rect 1135 37 1151 71
rect 1219 37 1235 71
rect 1293 37 1309 71
rect 1377 37 1393 71
rect 1451 37 1467 71
rect 1535 37 1551 71
rect 1609 37 1625 71
rect 1693 37 1709 71
rect 1767 37 1783 71
rect 1851 37 1867 71
rect 1925 37 1941 71
rect 2009 37 2025 71
rect 2083 37 2099 71
rect 2167 37 2183 71
rect -2183 -71 -2167 -37
rect -2099 -71 -2083 -37
rect -2025 -71 -2009 -37
rect -1941 -71 -1925 -37
rect -1867 -71 -1851 -37
rect -1783 -71 -1767 -37
rect -1709 -71 -1693 -37
rect -1625 -71 -1609 -37
rect -1551 -71 -1535 -37
rect -1467 -71 -1451 -37
rect -1393 -71 -1377 -37
rect -1309 -71 -1293 -37
rect -1235 -71 -1219 -37
rect -1151 -71 -1135 -37
rect -1077 -71 -1061 -37
rect -993 -71 -977 -37
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 977 -71 993 -37
rect 1061 -71 1077 -37
rect 1135 -71 1151 -37
rect 1219 -71 1235 -37
rect 1293 -71 1309 -37
rect 1377 -71 1393 -37
rect 1451 -71 1467 -37
rect 1535 -71 1551 -37
rect 1609 -71 1625 -37
rect 1693 -71 1709 -37
rect 1767 -71 1783 -37
rect 1851 -71 1867 -37
rect 1925 -71 1941 -37
rect 2009 -71 2025 -37
rect 2083 -71 2099 -37
rect 2167 -71 2183 -37
rect -2229 -121 -2195 -105
rect -2229 -1113 -2195 -1097
rect -2071 -121 -2037 -105
rect -2071 -1113 -2037 -1097
rect -1913 -121 -1879 -105
rect -1913 -1113 -1879 -1097
rect -1755 -121 -1721 -105
rect -1755 -1113 -1721 -1097
rect -1597 -121 -1563 -105
rect -1597 -1113 -1563 -1097
rect -1439 -121 -1405 -105
rect -1439 -1113 -1405 -1097
rect -1281 -121 -1247 -105
rect -1281 -1113 -1247 -1097
rect -1123 -121 -1089 -105
rect -1123 -1113 -1089 -1097
rect -965 -121 -931 -105
rect -965 -1113 -931 -1097
rect -807 -121 -773 -105
rect -807 -1113 -773 -1097
rect -649 -121 -615 -105
rect -649 -1113 -615 -1097
rect -491 -121 -457 -105
rect -491 -1113 -457 -1097
rect -333 -121 -299 -105
rect -333 -1113 -299 -1097
rect -175 -121 -141 -105
rect -175 -1113 -141 -1097
rect -17 -121 17 -105
rect -17 -1113 17 -1097
rect 141 -121 175 -105
rect 141 -1113 175 -1097
rect 299 -121 333 -105
rect 299 -1113 333 -1097
rect 457 -121 491 -105
rect 457 -1113 491 -1097
rect 615 -121 649 -105
rect 615 -1113 649 -1097
rect 773 -121 807 -105
rect 773 -1113 807 -1097
rect 931 -121 965 -105
rect 931 -1113 965 -1097
rect 1089 -121 1123 -105
rect 1089 -1113 1123 -1097
rect 1247 -121 1281 -105
rect 1247 -1113 1281 -1097
rect 1405 -121 1439 -105
rect 1405 -1113 1439 -1097
rect 1563 -121 1597 -105
rect 1563 -1113 1597 -1097
rect 1721 -121 1755 -105
rect 1721 -1113 1755 -1097
rect 1879 -121 1913 -105
rect 1879 -1113 1913 -1097
rect 2037 -121 2071 -105
rect 2037 -1113 2071 -1097
rect 2195 -121 2229 -105
rect 2195 -1113 2229 -1097
rect -2183 -1181 -2167 -1147
rect -2099 -1181 -2083 -1147
rect -2025 -1181 -2009 -1147
rect -1941 -1181 -1925 -1147
rect -1867 -1181 -1851 -1147
rect -1783 -1181 -1767 -1147
rect -1709 -1181 -1693 -1147
rect -1625 -1181 -1609 -1147
rect -1551 -1181 -1535 -1147
rect -1467 -1181 -1451 -1147
rect -1393 -1181 -1377 -1147
rect -1309 -1181 -1293 -1147
rect -1235 -1181 -1219 -1147
rect -1151 -1181 -1135 -1147
rect -1077 -1181 -1061 -1147
rect -993 -1181 -977 -1147
rect -919 -1181 -903 -1147
rect -835 -1181 -819 -1147
rect -761 -1181 -745 -1147
rect -677 -1181 -661 -1147
rect -603 -1181 -587 -1147
rect -519 -1181 -503 -1147
rect -445 -1181 -429 -1147
rect -361 -1181 -345 -1147
rect -287 -1181 -271 -1147
rect -203 -1181 -187 -1147
rect -129 -1181 -113 -1147
rect -45 -1181 -29 -1147
rect 29 -1181 45 -1147
rect 113 -1181 129 -1147
rect 187 -1181 203 -1147
rect 271 -1181 287 -1147
rect 345 -1181 361 -1147
rect 429 -1181 445 -1147
rect 503 -1181 519 -1147
rect 587 -1181 603 -1147
rect 661 -1181 677 -1147
rect 745 -1181 761 -1147
rect 819 -1181 835 -1147
rect 903 -1181 919 -1147
rect 977 -1181 993 -1147
rect 1061 -1181 1077 -1147
rect 1135 -1181 1151 -1147
rect 1219 -1181 1235 -1147
rect 1293 -1181 1309 -1147
rect 1377 -1181 1393 -1147
rect 1451 -1181 1467 -1147
rect 1535 -1181 1551 -1147
rect 1609 -1181 1625 -1147
rect 1693 -1181 1709 -1147
rect 1767 -1181 1783 -1147
rect 1851 -1181 1867 -1147
rect 1925 -1181 1941 -1147
rect 2009 -1181 2025 -1147
rect 2083 -1181 2099 -1147
rect 2167 -1181 2183 -1147
rect -2363 -1285 -2329 -1223
rect 2329 -1285 2363 -1223
rect -2363 -1319 -2267 -1285
rect 2267 -1319 2363 -1285
<< viali >>
rect -2167 1147 -2099 1181
rect -2009 1147 -1941 1181
rect -1851 1147 -1783 1181
rect -1693 1147 -1625 1181
rect -1535 1147 -1467 1181
rect -1377 1147 -1309 1181
rect -1219 1147 -1151 1181
rect -1061 1147 -993 1181
rect -903 1147 -835 1181
rect -745 1147 -677 1181
rect -587 1147 -519 1181
rect -429 1147 -361 1181
rect -271 1147 -203 1181
rect -113 1147 -45 1181
rect 45 1147 113 1181
rect 203 1147 271 1181
rect 361 1147 429 1181
rect 519 1147 587 1181
rect 677 1147 745 1181
rect 835 1147 903 1181
rect 993 1147 1061 1181
rect 1151 1147 1219 1181
rect 1309 1147 1377 1181
rect 1467 1147 1535 1181
rect 1625 1147 1693 1181
rect 1783 1147 1851 1181
rect 1941 1147 2009 1181
rect 2099 1147 2167 1181
rect -2229 121 -2195 1097
rect -2071 121 -2037 1097
rect -1913 121 -1879 1097
rect -1755 121 -1721 1097
rect -1597 121 -1563 1097
rect -1439 121 -1405 1097
rect -1281 121 -1247 1097
rect -1123 121 -1089 1097
rect -965 121 -931 1097
rect -807 121 -773 1097
rect -649 121 -615 1097
rect -491 121 -457 1097
rect -333 121 -299 1097
rect -175 121 -141 1097
rect -17 121 17 1097
rect 141 121 175 1097
rect 299 121 333 1097
rect 457 121 491 1097
rect 615 121 649 1097
rect 773 121 807 1097
rect 931 121 965 1097
rect 1089 121 1123 1097
rect 1247 121 1281 1097
rect 1405 121 1439 1097
rect 1563 121 1597 1097
rect 1721 121 1755 1097
rect 1879 121 1913 1097
rect 2037 121 2071 1097
rect 2195 121 2229 1097
rect -2167 37 -2099 71
rect -2009 37 -1941 71
rect -1851 37 -1783 71
rect -1693 37 -1625 71
rect -1535 37 -1467 71
rect -1377 37 -1309 71
rect -1219 37 -1151 71
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect 1151 37 1219 71
rect 1309 37 1377 71
rect 1467 37 1535 71
rect 1625 37 1693 71
rect 1783 37 1851 71
rect 1941 37 2009 71
rect 2099 37 2167 71
rect -2167 -71 -2099 -37
rect -2009 -71 -1941 -37
rect -1851 -71 -1783 -37
rect -1693 -71 -1625 -37
rect -1535 -71 -1467 -37
rect -1377 -71 -1309 -37
rect -1219 -71 -1151 -37
rect -1061 -71 -993 -37
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect 993 -71 1061 -37
rect 1151 -71 1219 -37
rect 1309 -71 1377 -37
rect 1467 -71 1535 -37
rect 1625 -71 1693 -37
rect 1783 -71 1851 -37
rect 1941 -71 2009 -37
rect 2099 -71 2167 -37
rect -2229 -1097 -2195 -121
rect -2071 -1097 -2037 -121
rect -1913 -1097 -1879 -121
rect -1755 -1097 -1721 -121
rect -1597 -1097 -1563 -121
rect -1439 -1097 -1405 -121
rect -1281 -1097 -1247 -121
rect -1123 -1097 -1089 -121
rect -965 -1097 -931 -121
rect -807 -1097 -773 -121
rect -649 -1097 -615 -121
rect -491 -1097 -457 -121
rect -333 -1097 -299 -121
rect -175 -1097 -141 -121
rect -17 -1097 17 -121
rect 141 -1097 175 -121
rect 299 -1097 333 -121
rect 457 -1097 491 -121
rect 615 -1097 649 -121
rect 773 -1097 807 -121
rect 931 -1097 965 -121
rect 1089 -1097 1123 -121
rect 1247 -1097 1281 -121
rect 1405 -1097 1439 -121
rect 1563 -1097 1597 -121
rect 1721 -1097 1755 -121
rect 1879 -1097 1913 -121
rect 2037 -1097 2071 -121
rect 2195 -1097 2229 -121
rect -2167 -1181 -2099 -1147
rect -2009 -1181 -1941 -1147
rect -1851 -1181 -1783 -1147
rect -1693 -1181 -1625 -1147
rect -1535 -1181 -1467 -1147
rect -1377 -1181 -1309 -1147
rect -1219 -1181 -1151 -1147
rect -1061 -1181 -993 -1147
rect -903 -1181 -835 -1147
rect -745 -1181 -677 -1147
rect -587 -1181 -519 -1147
rect -429 -1181 -361 -1147
rect -271 -1181 -203 -1147
rect -113 -1181 -45 -1147
rect 45 -1181 113 -1147
rect 203 -1181 271 -1147
rect 361 -1181 429 -1147
rect 519 -1181 587 -1147
rect 677 -1181 745 -1147
rect 835 -1181 903 -1147
rect 993 -1181 1061 -1147
rect 1151 -1181 1219 -1147
rect 1309 -1181 1377 -1147
rect 1467 -1181 1535 -1147
rect 1625 -1181 1693 -1147
rect 1783 -1181 1851 -1147
rect 1941 -1181 2009 -1147
rect 2099 -1181 2167 -1147
<< metal1 >>
rect -2179 1181 -2087 1187
rect -2179 1147 -2167 1181
rect -2099 1147 -2087 1181
rect -2179 1141 -2087 1147
rect -2021 1181 -1929 1187
rect -2021 1147 -2009 1181
rect -1941 1147 -1929 1181
rect -2021 1141 -1929 1147
rect -1863 1181 -1771 1187
rect -1863 1147 -1851 1181
rect -1783 1147 -1771 1181
rect -1863 1141 -1771 1147
rect -1705 1181 -1613 1187
rect -1705 1147 -1693 1181
rect -1625 1147 -1613 1181
rect -1705 1141 -1613 1147
rect -1547 1181 -1455 1187
rect -1547 1147 -1535 1181
rect -1467 1147 -1455 1181
rect -1547 1141 -1455 1147
rect -1389 1181 -1297 1187
rect -1389 1147 -1377 1181
rect -1309 1147 -1297 1181
rect -1389 1141 -1297 1147
rect -1231 1181 -1139 1187
rect -1231 1147 -1219 1181
rect -1151 1147 -1139 1181
rect -1231 1141 -1139 1147
rect -1073 1181 -981 1187
rect -1073 1147 -1061 1181
rect -993 1147 -981 1181
rect -1073 1141 -981 1147
rect -915 1181 -823 1187
rect -915 1147 -903 1181
rect -835 1147 -823 1181
rect -915 1141 -823 1147
rect -757 1181 -665 1187
rect -757 1147 -745 1181
rect -677 1147 -665 1181
rect -757 1141 -665 1147
rect -599 1181 -507 1187
rect -599 1147 -587 1181
rect -519 1147 -507 1181
rect -599 1141 -507 1147
rect -441 1181 -349 1187
rect -441 1147 -429 1181
rect -361 1147 -349 1181
rect -441 1141 -349 1147
rect -283 1181 -191 1187
rect -283 1147 -271 1181
rect -203 1147 -191 1181
rect -283 1141 -191 1147
rect -125 1181 -33 1187
rect -125 1147 -113 1181
rect -45 1147 -33 1181
rect -125 1141 -33 1147
rect 33 1181 125 1187
rect 33 1147 45 1181
rect 113 1147 125 1181
rect 33 1141 125 1147
rect 191 1181 283 1187
rect 191 1147 203 1181
rect 271 1147 283 1181
rect 191 1141 283 1147
rect 349 1181 441 1187
rect 349 1147 361 1181
rect 429 1147 441 1181
rect 349 1141 441 1147
rect 507 1181 599 1187
rect 507 1147 519 1181
rect 587 1147 599 1181
rect 507 1141 599 1147
rect 665 1181 757 1187
rect 665 1147 677 1181
rect 745 1147 757 1181
rect 665 1141 757 1147
rect 823 1181 915 1187
rect 823 1147 835 1181
rect 903 1147 915 1181
rect 823 1141 915 1147
rect 981 1181 1073 1187
rect 981 1147 993 1181
rect 1061 1147 1073 1181
rect 981 1141 1073 1147
rect 1139 1181 1231 1187
rect 1139 1147 1151 1181
rect 1219 1147 1231 1181
rect 1139 1141 1231 1147
rect 1297 1181 1389 1187
rect 1297 1147 1309 1181
rect 1377 1147 1389 1181
rect 1297 1141 1389 1147
rect 1455 1181 1547 1187
rect 1455 1147 1467 1181
rect 1535 1147 1547 1181
rect 1455 1141 1547 1147
rect 1613 1181 1705 1187
rect 1613 1147 1625 1181
rect 1693 1147 1705 1181
rect 1613 1141 1705 1147
rect 1771 1181 1863 1187
rect 1771 1147 1783 1181
rect 1851 1147 1863 1181
rect 1771 1141 1863 1147
rect 1929 1181 2021 1187
rect 1929 1147 1941 1181
rect 2009 1147 2021 1181
rect 1929 1141 2021 1147
rect 2087 1181 2179 1187
rect 2087 1147 2099 1181
rect 2167 1147 2179 1181
rect 2087 1141 2179 1147
rect -2235 1097 -2189 1109
rect -2235 121 -2229 1097
rect -2195 121 -2189 1097
rect -2235 109 -2189 121
rect -2077 1097 -2031 1109
rect -2077 121 -2071 1097
rect -2037 121 -2031 1097
rect -2077 109 -2031 121
rect -1919 1097 -1873 1109
rect -1919 121 -1913 1097
rect -1879 121 -1873 1097
rect -1919 109 -1873 121
rect -1761 1097 -1715 1109
rect -1761 121 -1755 1097
rect -1721 121 -1715 1097
rect -1761 109 -1715 121
rect -1603 1097 -1557 1109
rect -1603 121 -1597 1097
rect -1563 121 -1557 1097
rect -1603 109 -1557 121
rect -1445 1097 -1399 1109
rect -1445 121 -1439 1097
rect -1405 121 -1399 1097
rect -1445 109 -1399 121
rect -1287 1097 -1241 1109
rect -1287 121 -1281 1097
rect -1247 121 -1241 1097
rect -1287 109 -1241 121
rect -1129 1097 -1083 1109
rect -1129 121 -1123 1097
rect -1089 121 -1083 1097
rect -1129 109 -1083 121
rect -971 1097 -925 1109
rect -971 121 -965 1097
rect -931 121 -925 1097
rect -971 109 -925 121
rect -813 1097 -767 1109
rect -813 121 -807 1097
rect -773 121 -767 1097
rect -813 109 -767 121
rect -655 1097 -609 1109
rect -655 121 -649 1097
rect -615 121 -609 1097
rect -655 109 -609 121
rect -497 1097 -451 1109
rect -497 121 -491 1097
rect -457 121 -451 1097
rect -497 109 -451 121
rect -339 1097 -293 1109
rect -339 121 -333 1097
rect -299 121 -293 1097
rect -339 109 -293 121
rect -181 1097 -135 1109
rect -181 121 -175 1097
rect -141 121 -135 1097
rect -181 109 -135 121
rect -23 1097 23 1109
rect -23 121 -17 1097
rect 17 121 23 1097
rect -23 109 23 121
rect 135 1097 181 1109
rect 135 121 141 1097
rect 175 121 181 1097
rect 135 109 181 121
rect 293 1097 339 1109
rect 293 121 299 1097
rect 333 121 339 1097
rect 293 109 339 121
rect 451 1097 497 1109
rect 451 121 457 1097
rect 491 121 497 1097
rect 451 109 497 121
rect 609 1097 655 1109
rect 609 121 615 1097
rect 649 121 655 1097
rect 609 109 655 121
rect 767 1097 813 1109
rect 767 121 773 1097
rect 807 121 813 1097
rect 767 109 813 121
rect 925 1097 971 1109
rect 925 121 931 1097
rect 965 121 971 1097
rect 925 109 971 121
rect 1083 1097 1129 1109
rect 1083 121 1089 1097
rect 1123 121 1129 1097
rect 1083 109 1129 121
rect 1241 1097 1287 1109
rect 1241 121 1247 1097
rect 1281 121 1287 1097
rect 1241 109 1287 121
rect 1399 1097 1445 1109
rect 1399 121 1405 1097
rect 1439 121 1445 1097
rect 1399 109 1445 121
rect 1557 1097 1603 1109
rect 1557 121 1563 1097
rect 1597 121 1603 1097
rect 1557 109 1603 121
rect 1715 1097 1761 1109
rect 1715 121 1721 1097
rect 1755 121 1761 1097
rect 1715 109 1761 121
rect 1873 1097 1919 1109
rect 1873 121 1879 1097
rect 1913 121 1919 1097
rect 1873 109 1919 121
rect 2031 1097 2077 1109
rect 2031 121 2037 1097
rect 2071 121 2077 1097
rect 2031 109 2077 121
rect 2189 1097 2235 1109
rect 2189 121 2195 1097
rect 2229 121 2235 1097
rect 2189 109 2235 121
rect -2179 71 -2087 77
rect -2179 37 -2167 71
rect -2099 37 -2087 71
rect -2179 31 -2087 37
rect -2021 71 -1929 77
rect -2021 37 -2009 71
rect -1941 37 -1929 71
rect -2021 31 -1929 37
rect -1863 71 -1771 77
rect -1863 37 -1851 71
rect -1783 37 -1771 71
rect -1863 31 -1771 37
rect -1705 71 -1613 77
rect -1705 37 -1693 71
rect -1625 37 -1613 71
rect -1705 31 -1613 37
rect -1547 71 -1455 77
rect -1547 37 -1535 71
rect -1467 37 -1455 71
rect -1547 31 -1455 37
rect -1389 71 -1297 77
rect -1389 37 -1377 71
rect -1309 37 -1297 71
rect -1389 31 -1297 37
rect -1231 71 -1139 77
rect -1231 37 -1219 71
rect -1151 37 -1139 71
rect -1231 31 -1139 37
rect -1073 71 -981 77
rect -1073 37 -1061 71
rect -993 37 -981 71
rect -1073 31 -981 37
rect -915 71 -823 77
rect -915 37 -903 71
rect -835 37 -823 71
rect -915 31 -823 37
rect -757 71 -665 77
rect -757 37 -745 71
rect -677 37 -665 71
rect -757 31 -665 37
rect -599 71 -507 77
rect -599 37 -587 71
rect -519 37 -507 71
rect -599 31 -507 37
rect -441 71 -349 77
rect -441 37 -429 71
rect -361 37 -349 71
rect -441 31 -349 37
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect 349 71 441 77
rect 349 37 361 71
rect 429 37 441 71
rect 349 31 441 37
rect 507 71 599 77
rect 507 37 519 71
rect 587 37 599 71
rect 507 31 599 37
rect 665 71 757 77
rect 665 37 677 71
rect 745 37 757 71
rect 665 31 757 37
rect 823 71 915 77
rect 823 37 835 71
rect 903 37 915 71
rect 823 31 915 37
rect 981 71 1073 77
rect 981 37 993 71
rect 1061 37 1073 71
rect 981 31 1073 37
rect 1139 71 1231 77
rect 1139 37 1151 71
rect 1219 37 1231 71
rect 1139 31 1231 37
rect 1297 71 1389 77
rect 1297 37 1309 71
rect 1377 37 1389 71
rect 1297 31 1389 37
rect 1455 71 1547 77
rect 1455 37 1467 71
rect 1535 37 1547 71
rect 1455 31 1547 37
rect 1613 71 1705 77
rect 1613 37 1625 71
rect 1693 37 1705 71
rect 1613 31 1705 37
rect 1771 71 1863 77
rect 1771 37 1783 71
rect 1851 37 1863 71
rect 1771 31 1863 37
rect 1929 71 2021 77
rect 1929 37 1941 71
rect 2009 37 2021 71
rect 1929 31 2021 37
rect 2087 71 2179 77
rect 2087 37 2099 71
rect 2167 37 2179 71
rect 2087 31 2179 37
rect -2179 -37 -2087 -31
rect -2179 -71 -2167 -37
rect -2099 -71 -2087 -37
rect -2179 -77 -2087 -71
rect -2021 -37 -1929 -31
rect -2021 -71 -2009 -37
rect -1941 -71 -1929 -37
rect -2021 -77 -1929 -71
rect -1863 -37 -1771 -31
rect -1863 -71 -1851 -37
rect -1783 -71 -1771 -37
rect -1863 -77 -1771 -71
rect -1705 -37 -1613 -31
rect -1705 -71 -1693 -37
rect -1625 -71 -1613 -37
rect -1705 -77 -1613 -71
rect -1547 -37 -1455 -31
rect -1547 -71 -1535 -37
rect -1467 -71 -1455 -37
rect -1547 -77 -1455 -71
rect -1389 -37 -1297 -31
rect -1389 -71 -1377 -37
rect -1309 -71 -1297 -37
rect -1389 -77 -1297 -71
rect -1231 -37 -1139 -31
rect -1231 -71 -1219 -37
rect -1151 -71 -1139 -37
rect -1231 -77 -1139 -71
rect -1073 -37 -981 -31
rect -1073 -71 -1061 -37
rect -993 -71 -981 -37
rect -1073 -77 -981 -71
rect -915 -37 -823 -31
rect -915 -71 -903 -37
rect -835 -71 -823 -37
rect -915 -77 -823 -71
rect -757 -37 -665 -31
rect -757 -71 -745 -37
rect -677 -71 -665 -37
rect -757 -77 -665 -71
rect -599 -37 -507 -31
rect -599 -71 -587 -37
rect -519 -71 -507 -37
rect -599 -77 -507 -71
rect -441 -37 -349 -31
rect -441 -71 -429 -37
rect -361 -71 -349 -37
rect -441 -77 -349 -71
rect -283 -37 -191 -31
rect -283 -71 -271 -37
rect -203 -71 -191 -37
rect -283 -77 -191 -71
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect 191 -37 283 -31
rect 191 -71 203 -37
rect 271 -71 283 -37
rect 191 -77 283 -71
rect 349 -37 441 -31
rect 349 -71 361 -37
rect 429 -71 441 -37
rect 349 -77 441 -71
rect 507 -37 599 -31
rect 507 -71 519 -37
rect 587 -71 599 -37
rect 507 -77 599 -71
rect 665 -37 757 -31
rect 665 -71 677 -37
rect 745 -71 757 -37
rect 665 -77 757 -71
rect 823 -37 915 -31
rect 823 -71 835 -37
rect 903 -71 915 -37
rect 823 -77 915 -71
rect 981 -37 1073 -31
rect 981 -71 993 -37
rect 1061 -71 1073 -37
rect 981 -77 1073 -71
rect 1139 -37 1231 -31
rect 1139 -71 1151 -37
rect 1219 -71 1231 -37
rect 1139 -77 1231 -71
rect 1297 -37 1389 -31
rect 1297 -71 1309 -37
rect 1377 -71 1389 -37
rect 1297 -77 1389 -71
rect 1455 -37 1547 -31
rect 1455 -71 1467 -37
rect 1535 -71 1547 -37
rect 1455 -77 1547 -71
rect 1613 -37 1705 -31
rect 1613 -71 1625 -37
rect 1693 -71 1705 -37
rect 1613 -77 1705 -71
rect 1771 -37 1863 -31
rect 1771 -71 1783 -37
rect 1851 -71 1863 -37
rect 1771 -77 1863 -71
rect 1929 -37 2021 -31
rect 1929 -71 1941 -37
rect 2009 -71 2021 -37
rect 1929 -77 2021 -71
rect 2087 -37 2179 -31
rect 2087 -71 2099 -37
rect 2167 -71 2179 -37
rect 2087 -77 2179 -71
rect -2235 -121 -2189 -109
rect -2235 -1097 -2229 -121
rect -2195 -1097 -2189 -121
rect -2235 -1109 -2189 -1097
rect -2077 -121 -2031 -109
rect -2077 -1097 -2071 -121
rect -2037 -1097 -2031 -121
rect -2077 -1109 -2031 -1097
rect -1919 -121 -1873 -109
rect -1919 -1097 -1913 -121
rect -1879 -1097 -1873 -121
rect -1919 -1109 -1873 -1097
rect -1761 -121 -1715 -109
rect -1761 -1097 -1755 -121
rect -1721 -1097 -1715 -121
rect -1761 -1109 -1715 -1097
rect -1603 -121 -1557 -109
rect -1603 -1097 -1597 -121
rect -1563 -1097 -1557 -121
rect -1603 -1109 -1557 -1097
rect -1445 -121 -1399 -109
rect -1445 -1097 -1439 -121
rect -1405 -1097 -1399 -121
rect -1445 -1109 -1399 -1097
rect -1287 -121 -1241 -109
rect -1287 -1097 -1281 -121
rect -1247 -1097 -1241 -121
rect -1287 -1109 -1241 -1097
rect -1129 -121 -1083 -109
rect -1129 -1097 -1123 -121
rect -1089 -1097 -1083 -121
rect -1129 -1109 -1083 -1097
rect -971 -121 -925 -109
rect -971 -1097 -965 -121
rect -931 -1097 -925 -121
rect -971 -1109 -925 -1097
rect -813 -121 -767 -109
rect -813 -1097 -807 -121
rect -773 -1097 -767 -121
rect -813 -1109 -767 -1097
rect -655 -121 -609 -109
rect -655 -1097 -649 -121
rect -615 -1097 -609 -121
rect -655 -1109 -609 -1097
rect -497 -121 -451 -109
rect -497 -1097 -491 -121
rect -457 -1097 -451 -121
rect -497 -1109 -451 -1097
rect -339 -121 -293 -109
rect -339 -1097 -333 -121
rect -299 -1097 -293 -121
rect -339 -1109 -293 -1097
rect -181 -121 -135 -109
rect -181 -1097 -175 -121
rect -141 -1097 -135 -121
rect -181 -1109 -135 -1097
rect -23 -121 23 -109
rect -23 -1097 -17 -121
rect 17 -1097 23 -121
rect -23 -1109 23 -1097
rect 135 -121 181 -109
rect 135 -1097 141 -121
rect 175 -1097 181 -121
rect 135 -1109 181 -1097
rect 293 -121 339 -109
rect 293 -1097 299 -121
rect 333 -1097 339 -121
rect 293 -1109 339 -1097
rect 451 -121 497 -109
rect 451 -1097 457 -121
rect 491 -1097 497 -121
rect 451 -1109 497 -1097
rect 609 -121 655 -109
rect 609 -1097 615 -121
rect 649 -1097 655 -121
rect 609 -1109 655 -1097
rect 767 -121 813 -109
rect 767 -1097 773 -121
rect 807 -1097 813 -121
rect 767 -1109 813 -1097
rect 925 -121 971 -109
rect 925 -1097 931 -121
rect 965 -1097 971 -121
rect 925 -1109 971 -1097
rect 1083 -121 1129 -109
rect 1083 -1097 1089 -121
rect 1123 -1097 1129 -121
rect 1083 -1109 1129 -1097
rect 1241 -121 1287 -109
rect 1241 -1097 1247 -121
rect 1281 -1097 1287 -121
rect 1241 -1109 1287 -1097
rect 1399 -121 1445 -109
rect 1399 -1097 1405 -121
rect 1439 -1097 1445 -121
rect 1399 -1109 1445 -1097
rect 1557 -121 1603 -109
rect 1557 -1097 1563 -121
rect 1597 -1097 1603 -121
rect 1557 -1109 1603 -1097
rect 1715 -121 1761 -109
rect 1715 -1097 1721 -121
rect 1755 -1097 1761 -121
rect 1715 -1109 1761 -1097
rect 1873 -121 1919 -109
rect 1873 -1097 1879 -121
rect 1913 -1097 1919 -121
rect 1873 -1109 1919 -1097
rect 2031 -121 2077 -109
rect 2031 -1097 2037 -121
rect 2071 -1097 2077 -121
rect 2031 -1109 2077 -1097
rect 2189 -121 2235 -109
rect 2189 -1097 2195 -121
rect 2229 -1097 2235 -121
rect 2189 -1109 2235 -1097
rect -2179 -1147 -2087 -1141
rect -2179 -1181 -2167 -1147
rect -2099 -1181 -2087 -1147
rect -2179 -1187 -2087 -1181
rect -2021 -1147 -1929 -1141
rect -2021 -1181 -2009 -1147
rect -1941 -1181 -1929 -1147
rect -2021 -1187 -1929 -1181
rect -1863 -1147 -1771 -1141
rect -1863 -1181 -1851 -1147
rect -1783 -1181 -1771 -1147
rect -1863 -1187 -1771 -1181
rect -1705 -1147 -1613 -1141
rect -1705 -1181 -1693 -1147
rect -1625 -1181 -1613 -1147
rect -1705 -1187 -1613 -1181
rect -1547 -1147 -1455 -1141
rect -1547 -1181 -1535 -1147
rect -1467 -1181 -1455 -1147
rect -1547 -1187 -1455 -1181
rect -1389 -1147 -1297 -1141
rect -1389 -1181 -1377 -1147
rect -1309 -1181 -1297 -1147
rect -1389 -1187 -1297 -1181
rect -1231 -1147 -1139 -1141
rect -1231 -1181 -1219 -1147
rect -1151 -1181 -1139 -1147
rect -1231 -1187 -1139 -1181
rect -1073 -1147 -981 -1141
rect -1073 -1181 -1061 -1147
rect -993 -1181 -981 -1147
rect -1073 -1187 -981 -1181
rect -915 -1147 -823 -1141
rect -915 -1181 -903 -1147
rect -835 -1181 -823 -1147
rect -915 -1187 -823 -1181
rect -757 -1147 -665 -1141
rect -757 -1181 -745 -1147
rect -677 -1181 -665 -1147
rect -757 -1187 -665 -1181
rect -599 -1147 -507 -1141
rect -599 -1181 -587 -1147
rect -519 -1181 -507 -1147
rect -599 -1187 -507 -1181
rect -441 -1147 -349 -1141
rect -441 -1181 -429 -1147
rect -361 -1181 -349 -1147
rect -441 -1187 -349 -1181
rect -283 -1147 -191 -1141
rect -283 -1181 -271 -1147
rect -203 -1181 -191 -1147
rect -283 -1187 -191 -1181
rect -125 -1147 -33 -1141
rect -125 -1181 -113 -1147
rect -45 -1181 -33 -1147
rect -125 -1187 -33 -1181
rect 33 -1147 125 -1141
rect 33 -1181 45 -1147
rect 113 -1181 125 -1147
rect 33 -1187 125 -1181
rect 191 -1147 283 -1141
rect 191 -1181 203 -1147
rect 271 -1181 283 -1147
rect 191 -1187 283 -1181
rect 349 -1147 441 -1141
rect 349 -1181 361 -1147
rect 429 -1181 441 -1147
rect 349 -1187 441 -1181
rect 507 -1147 599 -1141
rect 507 -1181 519 -1147
rect 587 -1181 599 -1147
rect 507 -1187 599 -1181
rect 665 -1147 757 -1141
rect 665 -1181 677 -1147
rect 745 -1181 757 -1147
rect 665 -1187 757 -1181
rect 823 -1147 915 -1141
rect 823 -1181 835 -1147
rect 903 -1181 915 -1147
rect 823 -1187 915 -1181
rect 981 -1147 1073 -1141
rect 981 -1181 993 -1147
rect 1061 -1181 1073 -1147
rect 981 -1187 1073 -1181
rect 1139 -1147 1231 -1141
rect 1139 -1181 1151 -1147
rect 1219 -1181 1231 -1147
rect 1139 -1187 1231 -1181
rect 1297 -1147 1389 -1141
rect 1297 -1181 1309 -1147
rect 1377 -1181 1389 -1147
rect 1297 -1187 1389 -1181
rect 1455 -1147 1547 -1141
rect 1455 -1181 1467 -1147
rect 1535 -1181 1547 -1147
rect 1455 -1187 1547 -1181
rect 1613 -1147 1705 -1141
rect 1613 -1181 1625 -1147
rect 1693 -1181 1705 -1147
rect 1613 -1187 1705 -1181
rect 1771 -1147 1863 -1141
rect 1771 -1181 1783 -1147
rect 1851 -1181 1863 -1147
rect 1771 -1187 1863 -1181
rect 1929 -1147 2021 -1141
rect 1929 -1181 1941 -1147
rect 2009 -1181 2021 -1147
rect 1929 -1187 2021 -1181
rect 2087 -1147 2179 -1141
rect 2087 -1181 2099 -1147
rect 2167 -1181 2179 -1147
rect 2087 -1187 2179 -1181
<< properties >>
string FIXED_BBOX -2346 -1302 2346 1302
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.50 m 2 nf 28 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
