/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_mosbius (
    input  wire       VGND,
    input  wire       VDPWR,    // 1.8v power supply
    input  wire       VAPWR,    // 3.3v power supply
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    inout  wire [7:0] ua,       // Analog pins, only ua[5:0] can be used
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

    tt_um_mosbius mosbius (
        .bus5(ua[4]),
	.bus4(ua[3]),
	.bus3(ua[2]),
	.bus2(ua[1]),
	.bus1(ua[0]),
	.ibias(ua[5]),
	.VAPWR(VAPWR),
	.VDPWR(VDPWR),
	.VGND(VGND),
	.clk(clk),
	.dat_in(ui_in[0]),
	.rst_n(ui_in[2]),
	.dat_out(uo_out[0]),
	.enable(ui_in[1])
        );

endmodule
