magic
tech sky130A
magscale 1 2
timestamp 1757730208
<< nwell >>
rect -1651 -1297 1651 1297
<< mvpmos >>
rect -1393 -1000 -1293 1000
rect -1235 -1000 -1135 1000
rect -1077 -1000 -977 1000
rect -919 -1000 -819 1000
rect -761 -1000 -661 1000
rect -603 -1000 -503 1000
rect -445 -1000 -345 1000
rect -287 -1000 -187 1000
rect -129 -1000 -29 1000
rect 29 -1000 129 1000
rect 187 -1000 287 1000
rect 345 -1000 445 1000
rect 503 -1000 603 1000
rect 661 -1000 761 1000
rect 819 -1000 919 1000
rect 977 -1000 1077 1000
rect 1135 -1000 1235 1000
rect 1293 -1000 1393 1000
<< mvpdiff >>
rect -1451 988 -1393 1000
rect -1451 -988 -1439 988
rect -1405 -988 -1393 988
rect -1451 -1000 -1393 -988
rect -1293 988 -1235 1000
rect -1293 -988 -1281 988
rect -1247 -988 -1235 988
rect -1293 -1000 -1235 -988
rect -1135 988 -1077 1000
rect -1135 -988 -1123 988
rect -1089 -988 -1077 988
rect -1135 -1000 -1077 -988
rect -977 988 -919 1000
rect -977 -988 -965 988
rect -931 -988 -919 988
rect -977 -1000 -919 -988
rect -819 988 -761 1000
rect -819 -988 -807 988
rect -773 -988 -761 988
rect -819 -1000 -761 -988
rect -661 988 -603 1000
rect -661 -988 -649 988
rect -615 -988 -603 988
rect -661 -1000 -603 -988
rect -503 988 -445 1000
rect -503 -988 -491 988
rect -457 -988 -445 988
rect -503 -1000 -445 -988
rect -345 988 -287 1000
rect -345 -988 -333 988
rect -299 -988 -287 988
rect -345 -1000 -287 -988
rect -187 988 -129 1000
rect -187 -988 -175 988
rect -141 -988 -129 988
rect -187 -1000 -129 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 129 988 187 1000
rect 129 -988 141 988
rect 175 -988 187 988
rect 129 -1000 187 -988
rect 287 988 345 1000
rect 287 -988 299 988
rect 333 -988 345 988
rect 287 -1000 345 -988
rect 445 988 503 1000
rect 445 -988 457 988
rect 491 -988 503 988
rect 445 -1000 503 -988
rect 603 988 661 1000
rect 603 -988 615 988
rect 649 -988 661 988
rect 603 -1000 661 -988
rect 761 988 819 1000
rect 761 -988 773 988
rect 807 -988 819 988
rect 761 -1000 819 -988
rect 919 988 977 1000
rect 919 -988 931 988
rect 965 -988 977 988
rect 919 -1000 977 -988
rect 1077 988 1135 1000
rect 1077 -988 1089 988
rect 1123 -988 1135 988
rect 1077 -1000 1135 -988
rect 1235 988 1293 1000
rect 1235 -988 1247 988
rect 1281 -988 1293 988
rect 1235 -1000 1293 -988
rect 1393 988 1451 1000
rect 1393 -988 1405 988
rect 1439 -988 1451 988
rect 1393 -1000 1451 -988
<< mvpdiffc >>
rect -1439 -988 -1405 988
rect -1281 -988 -1247 988
rect -1123 -988 -1089 988
rect -965 -988 -931 988
rect -807 -988 -773 988
rect -649 -988 -615 988
rect -491 -988 -457 988
rect -333 -988 -299 988
rect -175 -988 -141 988
rect -17 -988 17 988
rect 141 -988 175 988
rect 299 -988 333 988
rect 457 -988 491 988
rect 615 -988 649 988
rect 773 -988 807 988
rect 931 -988 965 988
rect 1089 -988 1123 988
rect 1247 -988 1281 988
rect 1405 -988 1439 988
<< mvnsubdiff >>
rect -1585 1219 1585 1231
rect -1585 1185 -1477 1219
rect 1477 1185 1585 1219
rect -1585 1173 1585 1185
rect -1585 1123 -1527 1173
rect -1585 -1123 -1573 1123
rect -1539 -1123 -1527 1123
rect 1527 1123 1585 1173
rect -1585 -1173 -1527 -1123
rect 1527 -1123 1539 1123
rect 1573 -1123 1585 1123
rect 1527 -1173 1585 -1123
rect -1585 -1185 1585 -1173
rect -1585 -1219 -1477 -1185
rect 1477 -1219 1585 -1185
rect -1585 -1231 1585 -1219
<< mvnsubdiffcont >>
rect -1477 1185 1477 1219
rect -1573 -1123 -1539 1123
rect 1539 -1123 1573 1123
rect -1477 -1219 1477 -1185
<< poly >>
rect -1393 1081 -1293 1097
rect -1393 1047 -1377 1081
rect -1309 1047 -1293 1081
rect -1393 1000 -1293 1047
rect -1235 1081 -1135 1097
rect -1235 1047 -1219 1081
rect -1151 1047 -1135 1081
rect -1235 1000 -1135 1047
rect -1077 1081 -977 1097
rect -1077 1047 -1061 1081
rect -993 1047 -977 1081
rect -1077 1000 -977 1047
rect -919 1081 -819 1097
rect -919 1047 -903 1081
rect -835 1047 -819 1081
rect -919 1000 -819 1047
rect -761 1081 -661 1097
rect -761 1047 -745 1081
rect -677 1047 -661 1081
rect -761 1000 -661 1047
rect -603 1081 -503 1097
rect -603 1047 -587 1081
rect -519 1047 -503 1081
rect -603 1000 -503 1047
rect -445 1081 -345 1097
rect -445 1047 -429 1081
rect -361 1047 -345 1081
rect -445 1000 -345 1047
rect -287 1081 -187 1097
rect -287 1047 -271 1081
rect -203 1047 -187 1081
rect -287 1000 -187 1047
rect -129 1081 -29 1097
rect -129 1047 -113 1081
rect -45 1047 -29 1081
rect -129 1000 -29 1047
rect 29 1081 129 1097
rect 29 1047 45 1081
rect 113 1047 129 1081
rect 29 1000 129 1047
rect 187 1081 287 1097
rect 187 1047 203 1081
rect 271 1047 287 1081
rect 187 1000 287 1047
rect 345 1081 445 1097
rect 345 1047 361 1081
rect 429 1047 445 1081
rect 345 1000 445 1047
rect 503 1081 603 1097
rect 503 1047 519 1081
rect 587 1047 603 1081
rect 503 1000 603 1047
rect 661 1081 761 1097
rect 661 1047 677 1081
rect 745 1047 761 1081
rect 661 1000 761 1047
rect 819 1081 919 1097
rect 819 1047 835 1081
rect 903 1047 919 1081
rect 819 1000 919 1047
rect 977 1081 1077 1097
rect 977 1047 993 1081
rect 1061 1047 1077 1081
rect 977 1000 1077 1047
rect 1135 1081 1235 1097
rect 1135 1047 1151 1081
rect 1219 1047 1235 1081
rect 1135 1000 1235 1047
rect 1293 1081 1393 1097
rect 1293 1047 1309 1081
rect 1377 1047 1393 1081
rect 1293 1000 1393 1047
rect -1393 -1047 -1293 -1000
rect -1393 -1081 -1377 -1047
rect -1309 -1081 -1293 -1047
rect -1393 -1097 -1293 -1081
rect -1235 -1047 -1135 -1000
rect -1235 -1081 -1219 -1047
rect -1151 -1081 -1135 -1047
rect -1235 -1097 -1135 -1081
rect -1077 -1047 -977 -1000
rect -1077 -1081 -1061 -1047
rect -993 -1081 -977 -1047
rect -1077 -1097 -977 -1081
rect -919 -1047 -819 -1000
rect -919 -1081 -903 -1047
rect -835 -1081 -819 -1047
rect -919 -1097 -819 -1081
rect -761 -1047 -661 -1000
rect -761 -1081 -745 -1047
rect -677 -1081 -661 -1047
rect -761 -1097 -661 -1081
rect -603 -1047 -503 -1000
rect -603 -1081 -587 -1047
rect -519 -1081 -503 -1047
rect -603 -1097 -503 -1081
rect -445 -1047 -345 -1000
rect -445 -1081 -429 -1047
rect -361 -1081 -345 -1047
rect -445 -1097 -345 -1081
rect -287 -1047 -187 -1000
rect -287 -1081 -271 -1047
rect -203 -1081 -187 -1047
rect -287 -1097 -187 -1081
rect -129 -1047 -29 -1000
rect -129 -1081 -113 -1047
rect -45 -1081 -29 -1047
rect -129 -1097 -29 -1081
rect 29 -1047 129 -1000
rect 29 -1081 45 -1047
rect 113 -1081 129 -1047
rect 29 -1097 129 -1081
rect 187 -1047 287 -1000
rect 187 -1081 203 -1047
rect 271 -1081 287 -1047
rect 187 -1097 287 -1081
rect 345 -1047 445 -1000
rect 345 -1081 361 -1047
rect 429 -1081 445 -1047
rect 345 -1097 445 -1081
rect 503 -1047 603 -1000
rect 503 -1081 519 -1047
rect 587 -1081 603 -1047
rect 503 -1097 603 -1081
rect 661 -1047 761 -1000
rect 661 -1081 677 -1047
rect 745 -1081 761 -1047
rect 661 -1097 761 -1081
rect 819 -1047 919 -1000
rect 819 -1081 835 -1047
rect 903 -1081 919 -1047
rect 819 -1097 919 -1081
rect 977 -1047 1077 -1000
rect 977 -1081 993 -1047
rect 1061 -1081 1077 -1047
rect 977 -1097 1077 -1081
rect 1135 -1047 1235 -1000
rect 1135 -1081 1151 -1047
rect 1219 -1081 1235 -1047
rect 1135 -1097 1235 -1081
rect 1293 -1047 1393 -1000
rect 1293 -1081 1309 -1047
rect 1377 -1081 1393 -1047
rect 1293 -1097 1393 -1081
<< polycont >>
rect -1377 1047 -1309 1081
rect -1219 1047 -1151 1081
rect -1061 1047 -993 1081
rect -903 1047 -835 1081
rect -745 1047 -677 1081
rect -587 1047 -519 1081
rect -429 1047 -361 1081
rect -271 1047 -203 1081
rect -113 1047 -45 1081
rect 45 1047 113 1081
rect 203 1047 271 1081
rect 361 1047 429 1081
rect 519 1047 587 1081
rect 677 1047 745 1081
rect 835 1047 903 1081
rect 993 1047 1061 1081
rect 1151 1047 1219 1081
rect 1309 1047 1377 1081
rect -1377 -1081 -1309 -1047
rect -1219 -1081 -1151 -1047
rect -1061 -1081 -993 -1047
rect -903 -1081 -835 -1047
rect -745 -1081 -677 -1047
rect -587 -1081 -519 -1047
rect -429 -1081 -361 -1047
rect -271 -1081 -203 -1047
rect -113 -1081 -45 -1047
rect 45 -1081 113 -1047
rect 203 -1081 271 -1047
rect 361 -1081 429 -1047
rect 519 -1081 587 -1047
rect 677 -1081 745 -1047
rect 835 -1081 903 -1047
rect 993 -1081 1061 -1047
rect 1151 -1081 1219 -1047
rect 1309 -1081 1377 -1047
<< locali >>
rect -1573 1185 -1477 1219
rect 1477 1185 1573 1219
rect -1573 1123 -1539 1185
rect 1539 1123 1573 1185
rect -1393 1047 -1377 1081
rect -1309 1047 -1293 1081
rect -1235 1047 -1219 1081
rect -1151 1047 -1135 1081
rect -1077 1047 -1061 1081
rect -993 1047 -977 1081
rect -919 1047 -903 1081
rect -835 1047 -819 1081
rect -761 1047 -745 1081
rect -677 1047 -661 1081
rect -603 1047 -587 1081
rect -519 1047 -503 1081
rect -445 1047 -429 1081
rect -361 1047 -345 1081
rect -287 1047 -271 1081
rect -203 1047 -187 1081
rect -129 1047 -113 1081
rect -45 1047 -29 1081
rect 29 1047 45 1081
rect 113 1047 129 1081
rect 187 1047 203 1081
rect 271 1047 287 1081
rect 345 1047 361 1081
rect 429 1047 445 1081
rect 503 1047 519 1081
rect 587 1047 603 1081
rect 661 1047 677 1081
rect 745 1047 761 1081
rect 819 1047 835 1081
rect 903 1047 919 1081
rect 977 1047 993 1081
rect 1061 1047 1077 1081
rect 1135 1047 1151 1081
rect 1219 1047 1235 1081
rect 1293 1047 1309 1081
rect 1377 1047 1393 1081
rect -1439 988 -1405 1004
rect -1439 -1004 -1405 -988
rect -1281 988 -1247 1004
rect -1281 -1004 -1247 -988
rect -1123 988 -1089 1004
rect -1123 -1004 -1089 -988
rect -965 988 -931 1004
rect -965 -1004 -931 -988
rect -807 988 -773 1004
rect -807 -1004 -773 -988
rect -649 988 -615 1004
rect -649 -1004 -615 -988
rect -491 988 -457 1004
rect -491 -1004 -457 -988
rect -333 988 -299 1004
rect -333 -1004 -299 -988
rect -175 988 -141 1004
rect -175 -1004 -141 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 141 988 175 1004
rect 141 -1004 175 -988
rect 299 988 333 1004
rect 299 -1004 333 -988
rect 457 988 491 1004
rect 457 -1004 491 -988
rect 615 988 649 1004
rect 615 -1004 649 -988
rect 773 988 807 1004
rect 773 -1004 807 -988
rect 931 988 965 1004
rect 931 -1004 965 -988
rect 1089 988 1123 1004
rect 1089 -1004 1123 -988
rect 1247 988 1281 1004
rect 1247 -1004 1281 -988
rect 1405 988 1439 1004
rect 1405 -1004 1439 -988
rect -1393 -1081 -1377 -1047
rect -1309 -1081 -1293 -1047
rect -1235 -1081 -1219 -1047
rect -1151 -1081 -1135 -1047
rect -1077 -1081 -1061 -1047
rect -993 -1081 -977 -1047
rect -919 -1081 -903 -1047
rect -835 -1081 -819 -1047
rect -761 -1081 -745 -1047
rect -677 -1081 -661 -1047
rect -603 -1081 -587 -1047
rect -519 -1081 -503 -1047
rect -445 -1081 -429 -1047
rect -361 -1081 -345 -1047
rect -287 -1081 -271 -1047
rect -203 -1081 -187 -1047
rect -129 -1081 -113 -1047
rect -45 -1081 -29 -1047
rect 29 -1081 45 -1047
rect 113 -1081 129 -1047
rect 187 -1081 203 -1047
rect 271 -1081 287 -1047
rect 345 -1081 361 -1047
rect 429 -1081 445 -1047
rect 503 -1081 519 -1047
rect 587 -1081 603 -1047
rect 661 -1081 677 -1047
rect 745 -1081 761 -1047
rect 819 -1081 835 -1047
rect 903 -1081 919 -1047
rect 977 -1081 993 -1047
rect 1061 -1081 1077 -1047
rect 1135 -1081 1151 -1047
rect 1219 -1081 1235 -1047
rect 1293 -1081 1309 -1047
rect 1377 -1081 1393 -1047
rect -1573 -1185 -1539 -1123
rect 1539 -1185 1573 -1123
rect -1573 -1219 -1477 -1185
rect 1477 -1219 1573 -1185
<< viali >>
rect -1377 1047 -1309 1081
rect -1219 1047 -1151 1081
rect -1061 1047 -993 1081
rect -903 1047 -835 1081
rect -745 1047 -677 1081
rect -587 1047 -519 1081
rect -429 1047 -361 1081
rect -271 1047 -203 1081
rect -113 1047 -45 1081
rect 45 1047 113 1081
rect 203 1047 271 1081
rect 361 1047 429 1081
rect 519 1047 587 1081
rect 677 1047 745 1081
rect 835 1047 903 1081
rect 993 1047 1061 1081
rect 1151 1047 1219 1081
rect 1309 1047 1377 1081
rect -1439 -988 -1405 988
rect -1281 -988 -1247 988
rect -1123 -988 -1089 988
rect -965 -988 -931 988
rect -807 -988 -773 988
rect -649 -988 -615 988
rect -491 -988 -457 988
rect -333 -988 -299 988
rect -175 -988 -141 988
rect -17 -988 17 988
rect 141 -988 175 988
rect 299 -988 333 988
rect 457 -988 491 988
rect 615 -988 649 988
rect 773 -988 807 988
rect 931 -988 965 988
rect 1089 -988 1123 988
rect 1247 -988 1281 988
rect 1405 -988 1439 988
rect -1377 -1081 -1309 -1047
rect -1219 -1081 -1151 -1047
rect -1061 -1081 -993 -1047
rect -903 -1081 -835 -1047
rect -745 -1081 -677 -1047
rect -587 -1081 -519 -1047
rect -429 -1081 -361 -1047
rect -271 -1081 -203 -1047
rect -113 -1081 -45 -1047
rect 45 -1081 113 -1047
rect 203 -1081 271 -1047
rect 361 -1081 429 -1047
rect 519 -1081 587 -1047
rect 677 -1081 745 -1047
rect 835 -1081 903 -1047
rect 993 -1081 1061 -1047
rect 1151 -1081 1219 -1047
rect 1309 -1081 1377 -1047
<< metal1 >>
rect -1389 1081 -1297 1087
rect -1389 1047 -1377 1081
rect -1309 1047 -1297 1081
rect -1389 1041 -1297 1047
rect -1231 1081 -1139 1087
rect -1231 1047 -1219 1081
rect -1151 1047 -1139 1081
rect -1231 1041 -1139 1047
rect -1073 1081 -981 1087
rect -1073 1047 -1061 1081
rect -993 1047 -981 1081
rect -1073 1041 -981 1047
rect -915 1081 -823 1087
rect -915 1047 -903 1081
rect -835 1047 -823 1081
rect -915 1041 -823 1047
rect -757 1081 -665 1087
rect -757 1047 -745 1081
rect -677 1047 -665 1081
rect -757 1041 -665 1047
rect -599 1081 -507 1087
rect -599 1047 -587 1081
rect -519 1047 -507 1081
rect -599 1041 -507 1047
rect -441 1081 -349 1087
rect -441 1047 -429 1081
rect -361 1047 -349 1081
rect -441 1041 -349 1047
rect -283 1081 -191 1087
rect -283 1047 -271 1081
rect -203 1047 -191 1081
rect -283 1041 -191 1047
rect -125 1081 -33 1087
rect -125 1047 -113 1081
rect -45 1047 -33 1081
rect -125 1041 -33 1047
rect 33 1081 125 1087
rect 33 1047 45 1081
rect 113 1047 125 1081
rect 33 1041 125 1047
rect 191 1081 283 1087
rect 191 1047 203 1081
rect 271 1047 283 1081
rect 191 1041 283 1047
rect 349 1081 441 1087
rect 349 1047 361 1081
rect 429 1047 441 1081
rect 349 1041 441 1047
rect 507 1081 599 1087
rect 507 1047 519 1081
rect 587 1047 599 1081
rect 507 1041 599 1047
rect 665 1081 757 1087
rect 665 1047 677 1081
rect 745 1047 757 1081
rect 665 1041 757 1047
rect 823 1081 915 1087
rect 823 1047 835 1081
rect 903 1047 915 1081
rect 823 1041 915 1047
rect 981 1081 1073 1087
rect 981 1047 993 1081
rect 1061 1047 1073 1081
rect 981 1041 1073 1047
rect 1139 1081 1231 1087
rect 1139 1047 1151 1081
rect 1219 1047 1231 1081
rect 1139 1041 1231 1047
rect 1297 1081 1389 1087
rect 1297 1047 1309 1081
rect 1377 1047 1389 1081
rect 1297 1041 1389 1047
rect -1445 988 -1399 1000
rect -1445 -988 -1439 988
rect -1405 -988 -1399 988
rect -1445 -1000 -1399 -988
rect -1287 988 -1241 1000
rect -1287 -988 -1281 988
rect -1247 -988 -1241 988
rect -1287 -1000 -1241 -988
rect -1129 988 -1083 1000
rect -1129 -988 -1123 988
rect -1089 -988 -1083 988
rect -1129 -1000 -1083 -988
rect -971 988 -925 1000
rect -971 -988 -965 988
rect -931 -988 -925 988
rect -971 -1000 -925 -988
rect -813 988 -767 1000
rect -813 -988 -807 988
rect -773 -988 -767 988
rect -813 -1000 -767 -988
rect -655 988 -609 1000
rect -655 -988 -649 988
rect -615 -988 -609 988
rect -655 -1000 -609 -988
rect -497 988 -451 1000
rect -497 -988 -491 988
rect -457 -988 -451 988
rect -497 -1000 -451 -988
rect -339 988 -293 1000
rect -339 -988 -333 988
rect -299 -988 -293 988
rect -339 -1000 -293 -988
rect -181 988 -135 1000
rect -181 -988 -175 988
rect -141 -988 -135 988
rect -181 -1000 -135 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 135 988 181 1000
rect 135 -988 141 988
rect 175 -988 181 988
rect 135 -1000 181 -988
rect 293 988 339 1000
rect 293 -988 299 988
rect 333 -988 339 988
rect 293 -1000 339 -988
rect 451 988 497 1000
rect 451 -988 457 988
rect 491 -988 497 988
rect 451 -1000 497 -988
rect 609 988 655 1000
rect 609 -988 615 988
rect 649 -988 655 988
rect 609 -1000 655 -988
rect 767 988 813 1000
rect 767 -988 773 988
rect 807 -988 813 988
rect 767 -1000 813 -988
rect 925 988 971 1000
rect 925 -988 931 988
rect 965 -988 971 988
rect 925 -1000 971 -988
rect 1083 988 1129 1000
rect 1083 -988 1089 988
rect 1123 -988 1129 988
rect 1083 -1000 1129 -988
rect 1241 988 1287 1000
rect 1241 -988 1247 988
rect 1281 -988 1287 988
rect 1241 -1000 1287 -988
rect 1399 988 1445 1000
rect 1399 -988 1405 988
rect 1439 -988 1445 988
rect 1399 -1000 1445 -988
rect -1389 -1047 -1297 -1041
rect -1389 -1081 -1377 -1047
rect -1309 -1081 -1297 -1047
rect -1389 -1087 -1297 -1081
rect -1231 -1047 -1139 -1041
rect -1231 -1081 -1219 -1047
rect -1151 -1081 -1139 -1047
rect -1231 -1087 -1139 -1081
rect -1073 -1047 -981 -1041
rect -1073 -1081 -1061 -1047
rect -993 -1081 -981 -1047
rect -1073 -1087 -981 -1081
rect -915 -1047 -823 -1041
rect -915 -1081 -903 -1047
rect -835 -1081 -823 -1047
rect -915 -1087 -823 -1081
rect -757 -1047 -665 -1041
rect -757 -1081 -745 -1047
rect -677 -1081 -665 -1047
rect -757 -1087 -665 -1081
rect -599 -1047 -507 -1041
rect -599 -1081 -587 -1047
rect -519 -1081 -507 -1047
rect -599 -1087 -507 -1081
rect -441 -1047 -349 -1041
rect -441 -1081 -429 -1047
rect -361 -1081 -349 -1047
rect -441 -1087 -349 -1081
rect -283 -1047 -191 -1041
rect -283 -1081 -271 -1047
rect -203 -1081 -191 -1047
rect -283 -1087 -191 -1081
rect -125 -1047 -33 -1041
rect -125 -1081 -113 -1047
rect -45 -1081 -33 -1047
rect -125 -1087 -33 -1081
rect 33 -1047 125 -1041
rect 33 -1081 45 -1047
rect 113 -1081 125 -1047
rect 33 -1087 125 -1081
rect 191 -1047 283 -1041
rect 191 -1081 203 -1047
rect 271 -1081 283 -1047
rect 191 -1087 283 -1081
rect 349 -1047 441 -1041
rect 349 -1081 361 -1047
rect 429 -1081 441 -1047
rect 349 -1087 441 -1081
rect 507 -1047 599 -1041
rect 507 -1081 519 -1047
rect 587 -1081 599 -1047
rect 507 -1087 599 -1081
rect 665 -1047 757 -1041
rect 665 -1081 677 -1047
rect 745 -1081 757 -1047
rect 665 -1087 757 -1081
rect 823 -1047 915 -1041
rect 823 -1081 835 -1047
rect 903 -1081 915 -1047
rect 823 -1087 915 -1081
rect 981 -1047 1073 -1041
rect 981 -1081 993 -1047
rect 1061 -1081 1073 -1047
rect 981 -1087 1073 -1081
rect 1139 -1047 1231 -1041
rect 1139 -1081 1151 -1047
rect 1219 -1081 1231 -1047
rect 1139 -1087 1231 -1081
rect 1297 -1047 1389 -1041
rect 1297 -1081 1309 -1047
rect 1377 -1081 1389 -1047
rect 1297 -1087 1389 -1081
<< properties >>
string FIXED_BBOX -1556 -1202 1556 1202
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10 l 0.5 m 1 nf 18 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
