magic
tech sky130A
magscale 1 2
timestamp 1757105855
<< nwell >>
rect -5127 -2651 5127 2651
<< mvpmos >>
rect -4869 1354 -4769 2354
rect -4711 1354 -4611 2354
rect -4553 1354 -4453 2354
rect -4395 1354 -4295 2354
rect -4237 1354 -4137 2354
rect -4079 1354 -3979 2354
rect -3921 1354 -3821 2354
rect -3763 1354 -3663 2354
rect -3605 1354 -3505 2354
rect -3447 1354 -3347 2354
rect -3289 1354 -3189 2354
rect -3131 1354 -3031 2354
rect -2973 1354 -2873 2354
rect -2815 1354 -2715 2354
rect -2657 1354 -2557 2354
rect -2499 1354 -2399 2354
rect -2341 1354 -2241 2354
rect -2183 1354 -2083 2354
rect -2025 1354 -1925 2354
rect -1867 1354 -1767 2354
rect -1709 1354 -1609 2354
rect -1551 1354 -1451 2354
rect -1393 1354 -1293 2354
rect -1235 1354 -1135 2354
rect -1077 1354 -977 2354
rect -919 1354 -819 2354
rect -761 1354 -661 2354
rect -603 1354 -503 2354
rect -445 1354 -345 2354
rect -287 1354 -187 2354
rect -129 1354 -29 2354
rect 29 1354 129 2354
rect 187 1354 287 2354
rect 345 1354 445 2354
rect 503 1354 603 2354
rect 661 1354 761 2354
rect 819 1354 919 2354
rect 977 1354 1077 2354
rect 1135 1354 1235 2354
rect 1293 1354 1393 2354
rect 1451 1354 1551 2354
rect 1609 1354 1709 2354
rect 1767 1354 1867 2354
rect 1925 1354 2025 2354
rect 2083 1354 2183 2354
rect 2241 1354 2341 2354
rect 2399 1354 2499 2354
rect 2557 1354 2657 2354
rect 2715 1354 2815 2354
rect 2873 1354 2973 2354
rect 3031 1354 3131 2354
rect 3189 1354 3289 2354
rect 3347 1354 3447 2354
rect 3505 1354 3605 2354
rect 3663 1354 3763 2354
rect 3821 1354 3921 2354
rect 3979 1354 4079 2354
rect 4137 1354 4237 2354
rect 4295 1354 4395 2354
rect 4453 1354 4553 2354
rect 4611 1354 4711 2354
rect 4769 1354 4869 2354
rect -4869 118 -4769 1118
rect -4711 118 -4611 1118
rect -4553 118 -4453 1118
rect -4395 118 -4295 1118
rect -4237 118 -4137 1118
rect -4079 118 -3979 1118
rect -3921 118 -3821 1118
rect -3763 118 -3663 1118
rect -3605 118 -3505 1118
rect -3447 118 -3347 1118
rect -3289 118 -3189 1118
rect -3131 118 -3031 1118
rect -2973 118 -2873 1118
rect -2815 118 -2715 1118
rect -2657 118 -2557 1118
rect -2499 118 -2399 1118
rect -2341 118 -2241 1118
rect -2183 118 -2083 1118
rect -2025 118 -1925 1118
rect -1867 118 -1767 1118
rect -1709 118 -1609 1118
rect -1551 118 -1451 1118
rect -1393 118 -1293 1118
rect -1235 118 -1135 1118
rect -1077 118 -977 1118
rect -919 118 -819 1118
rect -761 118 -661 1118
rect -603 118 -503 1118
rect -445 118 -345 1118
rect -287 118 -187 1118
rect -129 118 -29 1118
rect 29 118 129 1118
rect 187 118 287 1118
rect 345 118 445 1118
rect 503 118 603 1118
rect 661 118 761 1118
rect 819 118 919 1118
rect 977 118 1077 1118
rect 1135 118 1235 1118
rect 1293 118 1393 1118
rect 1451 118 1551 1118
rect 1609 118 1709 1118
rect 1767 118 1867 1118
rect 1925 118 2025 1118
rect 2083 118 2183 1118
rect 2241 118 2341 1118
rect 2399 118 2499 1118
rect 2557 118 2657 1118
rect 2715 118 2815 1118
rect 2873 118 2973 1118
rect 3031 118 3131 1118
rect 3189 118 3289 1118
rect 3347 118 3447 1118
rect 3505 118 3605 1118
rect 3663 118 3763 1118
rect 3821 118 3921 1118
rect 3979 118 4079 1118
rect 4137 118 4237 1118
rect 4295 118 4395 1118
rect 4453 118 4553 1118
rect 4611 118 4711 1118
rect 4769 118 4869 1118
rect -4869 -1118 -4769 -118
rect -4711 -1118 -4611 -118
rect -4553 -1118 -4453 -118
rect -4395 -1118 -4295 -118
rect -4237 -1118 -4137 -118
rect -4079 -1118 -3979 -118
rect -3921 -1118 -3821 -118
rect -3763 -1118 -3663 -118
rect -3605 -1118 -3505 -118
rect -3447 -1118 -3347 -118
rect -3289 -1118 -3189 -118
rect -3131 -1118 -3031 -118
rect -2973 -1118 -2873 -118
rect -2815 -1118 -2715 -118
rect -2657 -1118 -2557 -118
rect -2499 -1118 -2399 -118
rect -2341 -1118 -2241 -118
rect -2183 -1118 -2083 -118
rect -2025 -1118 -1925 -118
rect -1867 -1118 -1767 -118
rect -1709 -1118 -1609 -118
rect -1551 -1118 -1451 -118
rect -1393 -1118 -1293 -118
rect -1235 -1118 -1135 -118
rect -1077 -1118 -977 -118
rect -919 -1118 -819 -118
rect -761 -1118 -661 -118
rect -603 -1118 -503 -118
rect -445 -1118 -345 -118
rect -287 -1118 -187 -118
rect -129 -1118 -29 -118
rect 29 -1118 129 -118
rect 187 -1118 287 -118
rect 345 -1118 445 -118
rect 503 -1118 603 -118
rect 661 -1118 761 -118
rect 819 -1118 919 -118
rect 977 -1118 1077 -118
rect 1135 -1118 1235 -118
rect 1293 -1118 1393 -118
rect 1451 -1118 1551 -118
rect 1609 -1118 1709 -118
rect 1767 -1118 1867 -118
rect 1925 -1118 2025 -118
rect 2083 -1118 2183 -118
rect 2241 -1118 2341 -118
rect 2399 -1118 2499 -118
rect 2557 -1118 2657 -118
rect 2715 -1118 2815 -118
rect 2873 -1118 2973 -118
rect 3031 -1118 3131 -118
rect 3189 -1118 3289 -118
rect 3347 -1118 3447 -118
rect 3505 -1118 3605 -118
rect 3663 -1118 3763 -118
rect 3821 -1118 3921 -118
rect 3979 -1118 4079 -118
rect 4137 -1118 4237 -118
rect 4295 -1118 4395 -118
rect 4453 -1118 4553 -118
rect 4611 -1118 4711 -118
rect 4769 -1118 4869 -118
rect -4869 -2354 -4769 -1354
rect -4711 -2354 -4611 -1354
rect -4553 -2354 -4453 -1354
rect -4395 -2354 -4295 -1354
rect -4237 -2354 -4137 -1354
rect -4079 -2354 -3979 -1354
rect -3921 -2354 -3821 -1354
rect -3763 -2354 -3663 -1354
rect -3605 -2354 -3505 -1354
rect -3447 -2354 -3347 -1354
rect -3289 -2354 -3189 -1354
rect -3131 -2354 -3031 -1354
rect -2973 -2354 -2873 -1354
rect -2815 -2354 -2715 -1354
rect -2657 -2354 -2557 -1354
rect -2499 -2354 -2399 -1354
rect -2341 -2354 -2241 -1354
rect -2183 -2354 -2083 -1354
rect -2025 -2354 -1925 -1354
rect -1867 -2354 -1767 -1354
rect -1709 -2354 -1609 -1354
rect -1551 -2354 -1451 -1354
rect -1393 -2354 -1293 -1354
rect -1235 -2354 -1135 -1354
rect -1077 -2354 -977 -1354
rect -919 -2354 -819 -1354
rect -761 -2354 -661 -1354
rect -603 -2354 -503 -1354
rect -445 -2354 -345 -1354
rect -287 -2354 -187 -1354
rect -129 -2354 -29 -1354
rect 29 -2354 129 -1354
rect 187 -2354 287 -1354
rect 345 -2354 445 -1354
rect 503 -2354 603 -1354
rect 661 -2354 761 -1354
rect 819 -2354 919 -1354
rect 977 -2354 1077 -1354
rect 1135 -2354 1235 -1354
rect 1293 -2354 1393 -1354
rect 1451 -2354 1551 -1354
rect 1609 -2354 1709 -1354
rect 1767 -2354 1867 -1354
rect 1925 -2354 2025 -1354
rect 2083 -2354 2183 -1354
rect 2241 -2354 2341 -1354
rect 2399 -2354 2499 -1354
rect 2557 -2354 2657 -1354
rect 2715 -2354 2815 -1354
rect 2873 -2354 2973 -1354
rect 3031 -2354 3131 -1354
rect 3189 -2354 3289 -1354
rect 3347 -2354 3447 -1354
rect 3505 -2354 3605 -1354
rect 3663 -2354 3763 -1354
rect 3821 -2354 3921 -1354
rect 3979 -2354 4079 -1354
rect 4137 -2354 4237 -1354
rect 4295 -2354 4395 -1354
rect 4453 -2354 4553 -1354
rect 4611 -2354 4711 -1354
rect 4769 -2354 4869 -1354
<< mvpdiff >>
rect -4927 2342 -4869 2354
rect -4927 1366 -4915 2342
rect -4881 1366 -4869 2342
rect -4927 1354 -4869 1366
rect -4769 2342 -4711 2354
rect -4769 1366 -4757 2342
rect -4723 1366 -4711 2342
rect -4769 1354 -4711 1366
rect -4611 2342 -4553 2354
rect -4611 1366 -4599 2342
rect -4565 1366 -4553 2342
rect -4611 1354 -4553 1366
rect -4453 2342 -4395 2354
rect -4453 1366 -4441 2342
rect -4407 1366 -4395 2342
rect -4453 1354 -4395 1366
rect -4295 2342 -4237 2354
rect -4295 1366 -4283 2342
rect -4249 1366 -4237 2342
rect -4295 1354 -4237 1366
rect -4137 2342 -4079 2354
rect -4137 1366 -4125 2342
rect -4091 1366 -4079 2342
rect -4137 1354 -4079 1366
rect -3979 2342 -3921 2354
rect -3979 1366 -3967 2342
rect -3933 1366 -3921 2342
rect -3979 1354 -3921 1366
rect -3821 2342 -3763 2354
rect -3821 1366 -3809 2342
rect -3775 1366 -3763 2342
rect -3821 1354 -3763 1366
rect -3663 2342 -3605 2354
rect -3663 1366 -3651 2342
rect -3617 1366 -3605 2342
rect -3663 1354 -3605 1366
rect -3505 2342 -3447 2354
rect -3505 1366 -3493 2342
rect -3459 1366 -3447 2342
rect -3505 1354 -3447 1366
rect -3347 2342 -3289 2354
rect -3347 1366 -3335 2342
rect -3301 1366 -3289 2342
rect -3347 1354 -3289 1366
rect -3189 2342 -3131 2354
rect -3189 1366 -3177 2342
rect -3143 1366 -3131 2342
rect -3189 1354 -3131 1366
rect -3031 2342 -2973 2354
rect -3031 1366 -3019 2342
rect -2985 1366 -2973 2342
rect -3031 1354 -2973 1366
rect -2873 2342 -2815 2354
rect -2873 1366 -2861 2342
rect -2827 1366 -2815 2342
rect -2873 1354 -2815 1366
rect -2715 2342 -2657 2354
rect -2715 1366 -2703 2342
rect -2669 1366 -2657 2342
rect -2715 1354 -2657 1366
rect -2557 2342 -2499 2354
rect -2557 1366 -2545 2342
rect -2511 1366 -2499 2342
rect -2557 1354 -2499 1366
rect -2399 2342 -2341 2354
rect -2399 1366 -2387 2342
rect -2353 1366 -2341 2342
rect -2399 1354 -2341 1366
rect -2241 2342 -2183 2354
rect -2241 1366 -2229 2342
rect -2195 1366 -2183 2342
rect -2241 1354 -2183 1366
rect -2083 2342 -2025 2354
rect -2083 1366 -2071 2342
rect -2037 1366 -2025 2342
rect -2083 1354 -2025 1366
rect -1925 2342 -1867 2354
rect -1925 1366 -1913 2342
rect -1879 1366 -1867 2342
rect -1925 1354 -1867 1366
rect -1767 2342 -1709 2354
rect -1767 1366 -1755 2342
rect -1721 1366 -1709 2342
rect -1767 1354 -1709 1366
rect -1609 2342 -1551 2354
rect -1609 1366 -1597 2342
rect -1563 1366 -1551 2342
rect -1609 1354 -1551 1366
rect -1451 2342 -1393 2354
rect -1451 1366 -1439 2342
rect -1405 1366 -1393 2342
rect -1451 1354 -1393 1366
rect -1293 2342 -1235 2354
rect -1293 1366 -1281 2342
rect -1247 1366 -1235 2342
rect -1293 1354 -1235 1366
rect -1135 2342 -1077 2354
rect -1135 1366 -1123 2342
rect -1089 1366 -1077 2342
rect -1135 1354 -1077 1366
rect -977 2342 -919 2354
rect -977 1366 -965 2342
rect -931 1366 -919 2342
rect -977 1354 -919 1366
rect -819 2342 -761 2354
rect -819 1366 -807 2342
rect -773 1366 -761 2342
rect -819 1354 -761 1366
rect -661 2342 -603 2354
rect -661 1366 -649 2342
rect -615 1366 -603 2342
rect -661 1354 -603 1366
rect -503 2342 -445 2354
rect -503 1366 -491 2342
rect -457 1366 -445 2342
rect -503 1354 -445 1366
rect -345 2342 -287 2354
rect -345 1366 -333 2342
rect -299 1366 -287 2342
rect -345 1354 -287 1366
rect -187 2342 -129 2354
rect -187 1366 -175 2342
rect -141 1366 -129 2342
rect -187 1354 -129 1366
rect -29 2342 29 2354
rect -29 1366 -17 2342
rect 17 1366 29 2342
rect -29 1354 29 1366
rect 129 2342 187 2354
rect 129 1366 141 2342
rect 175 1366 187 2342
rect 129 1354 187 1366
rect 287 2342 345 2354
rect 287 1366 299 2342
rect 333 1366 345 2342
rect 287 1354 345 1366
rect 445 2342 503 2354
rect 445 1366 457 2342
rect 491 1366 503 2342
rect 445 1354 503 1366
rect 603 2342 661 2354
rect 603 1366 615 2342
rect 649 1366 661 2342
rect 603 1354 661 1366
rect 761 2342 819 2354
rect 761 1366 773 2342
rect 807 1366 819 2342
rect 761 1354 819 1366
rect 919 2342 977 2354
rect 919 1366 931 2342
rect 965 1366 977 2342
rect 919 1354 977 1366
rect 1077 2342 1135 2354
rect 1077 1366 1089 2342
rect 1123 1366 1135 2342
rect 1077 1354 1135 1366
rect 1235 2342 1293 2354
rect 1235 1366 1247 2342
rect 1281 1366 1293 2342
rect 1235 1354 1293 1366
rect 1393 2342 1451 2354
rect 1393 1366 1405 2342
rect 1439 1366 1451 2342
rect 1393 1354 1451 1366
rect 1551 2342 1609 2354
rect 1551 1366 1563 2342
rect 1597 1366 1609 2342
rect 1551 1354 1609 1366
rect 1709 2342 1767 2354
rect 1709 1366 1721 2342
rect 1755 1366 1767 2342
rect 1709 1354 1767 1366
rect 1867 2342 1925 2354
rect 1867 1366 1879 2342
rect 1913 1366 1925 2342
rect 1867 1354 1925 1366
rect 2025 2342 2083 2354
rect 2025 1366 2037 2342
rect 2071 1366 2083 2342
rect 2025 1354 2083 1366
rect 2183 2342 2241 2354
rect 2183 1366 2195 2342
rect 2229 1366 2241 2342
rect 2183 1354 2241 1366
rect 2341 2342 2399 2354
rect 2341 1366 2353 2342
rect 2387 1366 2399 2342
rect 2341 1354 2399 1366
rect 2499 2342 2557 2354
rect 2499 1366 2511 2342
rect 2545 1366 2557 2342
rect 2499 1354 2557 1366
rect 2657 2342 2715 2354
rect 2657 1366 2669 2342
rect 2703 1366 2715 2342
rect 2657 1354 2715 1366
rect 2815 2342 2873 2354
rect 2815 1366 2827 2342
rect 2861 1366 2873 2342
rect 2815 1354 2873 1366
rect 2973 2342 3031 2354
rect 2973 1366 2985 2342
rect 3019 1366 3031 2342
rect 2973 1354 3031 1366
rect 3131 2342 3189 2354
rect 3131 1366 3143 2342
rect 3177 1366 3189 2342
rect 3131 1354 3189 1366
rect 3289 2342 3347 2354
rect 3289 1366 3301 2342
rect 3335 1366 3347 2342
rect 3289 1354 3347 1366
rect 3447 2342 3505 2354
rect 3447 1366 3459 2342
rect 3493 1366 3505 2342
rect 3447 1354 3505 1366
rect 3605 2342 3663 2354
rect 3605 1366 3617 2342
rect 3651 1366 3663 2342
rect 3605 1354 3663 1366
rect 3763 2342 3821 2354
rect 3763 1366 3775 2342
rect 3809 1366 3821 2342
rect 3763 1354 3821 1366
rect 3921 2342 3979 2354
rect 3921 1366 3933 2342
rect 3967 1366 3979 2342
rect 3921 1354 3979 1366
rect 4079 2342 4137 2354
rect 4079 1366 4091 2342
rect 4125 1366 4137 2342
rect 4079 1354 4137 1366
rect 4237 2342 4295 2354
rect 4237 1366 4249 2342
rect 4283 1366 4295 2342
rect 4237 1354 4295 1366
rect 4395 2342 4453 2354
rect 4395 1366 4407 2342
rect 4441 1366 4453 2342
rect 4395 1354 4453 1366
rect 4553 2342 4611 2354
rect 4553 1366 4565 2342
rect 4599 1366 4611 2342
rect 4553 1354 4611 1366
rect 4711 2342 4769 2354
rect 4711 1366 4723 2342
rect 4757 1366 4769 2342
rect 4711 1354 4769 1366
rect 4869 2342 4927 2354
rect 4869 1366 4881 2342
rect 4915 1366 4927 2342
rect 4869 1354 4927 1366
rect -4927 1106 -4869 1118
rect -4927 130 -4915 1106
rect -4881 130 -4869 1106
rect -4927 118 -4869 130
rect -4769 1106 -4711 1118
rect -4769 130 -4757 1106
rect -4723 130 -4711 1106
rect -4769 118 -4711 130
rect -4611 1106 -4553 1118
rect -4611 130 -4599 1106
rect -4565 130 -4553 1106
rect -4611 118 -4553 130
rect -4453 1106 -4395 1118
rect -4453 130 -4441 1106
rect -4407 130 -4395 1106
rect -4453 118 -4395 130
rect -4295 1106 -4237 1118
rect -4295 130 -4283 1106
rect -4249 130 -4237 1106
rect -4295 118 -4237 130
rect -4137 1106 -4079 1118
rect -4137 130 -4125 1106
rect -4091 130 -4079 1106
rect -4137 118 -4079 130
rect -3979 1106 -3921 1118
rect -3979 130 -3967 1106
rect -3933 130 -3921 1106
rect -3979 118 -3921 130
rect -3821 1106 -3763 1118
rect -3821 130 -3809 1106
rect -3775 130 -3763 1106
rect -3821 118 -3763 130
rect -3663 1106 -3605 1118
rect -3663 130 -3651 1106
rect -3617 130 -3605 1106
rect -3663 118 -3605 130
rect -3505 1106 -3447 1118
rect -3505 130 -3493 1106
rect -3459 130 -3447 1106
rect -3505 118 -3447 130
rect -3347 1106 -3289 1118
rect -3347 130 -3335 1106
rect -3301 130 -3289 1106
rect -3347 118 -3289 130
rect -3189 1106 -3131 1118
rect -3189 130 -3177 1106
rect -3143 130 -3131 1106
rect -3189 118 -3131 130
rect -3031 1106 -2973 1118
rect -3031 130 -3019 1106
rect -2985 130 -2973 1106
rect -3031 118 -2973 130
rect -2873 1106 -2815 1118
rect -2873 130 -2861 1106
rect -2827 130 -2815 1106
rect -2873 118 -2815 130
rect -2715 1106 -2657 1118
rect -2715 130 -2703 1106
rect -2669 130 -2657 1106
rect -2715 118 -2657 130
rect -2557 1106 -2499 1118
rect -2557 130 -2545 1106
rect -2511 130 -2499 1106
rect -2557 118 -2499 130
rect -2399 1106 -2341 1118
rect -2399 130 -2387 1106
rect -2353 130 -2341 1106
rect -2399 118 -2341 130
rect -2241 1106 -2183 1118
rect -2241 130 -2229 1106
rect -2195 130 -2183 1106
rect -2241 118 -2183 130
rect -2083 1106 -2025 1118
rect -2083 130 -2071 1106
rect -2037 130 -2025 1106
rect -2083 118 -2025 130
rect -1925 1106 -1867 1118
rect -1925 130 -1913 1106
rect -1879 130 -1867 1106
rect -1925 118 -1867 130
rect -1767 1106 -1709 1118
rect -1767 130 -1755 1106
rect -1721 130 -1709 1106
rect -1767 118 -1709 130
rect -1609 1106 -1551 1118
rect -1609 130 -1597 1106
rect -1563 130 -1551 1106
rect -1609 118 -1551 130
rect -1451 1106 -1393 1118
rect -1451 130 -1439 1106
rect -1405 130 -1393 1106
rect -1451 118 -1393 130
rect -1293 1106 -1235 1118
rect -1293 130 -1281 1106
rect -1247 130 -1235 1106
rect -1293 118 -1235 130
rect -1135 1106 -1077 1118
rect -1135 130 -1123 1106
rect -1089 130 -1077 1106
rect -1135 118 -1077 130
rect -977 1106 -919 1118
rect -977 130 -965 1106
rect -931 130 -919 1106
rect -977 118 -919 130
rect -819 1106 -761 1118
rect -819 130 -807 1106
rect -773 130 -761 1106
rect -819 118 -761 130
rect -661 1106 -603 1118
rect -661 130 -649 1106
rect -615 130 -603 1106
rect -661 118 -603 130
rect -503 1106 -445 1118
rect -503 130 -491 1106
rect -457 130 -445 1106
rect -503 118 -445 130
rect -345 1106 -287 1118
rect -345 130 -333 1106
rect -299 130 -287 1106
rect -345 118 -287 130
rect -187 1106 -129 1118
rect -187 130 -175 1106
rect -141 130 -129 1106
rect -187 118 -129 130
rect -29 1106 29 1118
rect -29 130 -17 1106
rect 17 130 29 1106
rect -29 118 29 130
rect 129 1106 187 1118
rect 129 130 141 1106
rect 175 130 187 1106
rect 129 118 187 130
rect 287 1106 345 1118
rect 287 130 299 1106
rect 333 130 345 1106
rect 287 118 345 130
rect 445 1106 503 1118
rect 445 130 457 1106
rect 491 130 503 1106
rect 445 118 503 130
rect 603 1106 661 1118
rect 603 130 615 1106
rect 649 130 661 1106
rect 603 118 661 130
rect 761 1106 819 1118
rect 761 130 773 1106
rect 807 130 819 1106
rect 761 118 819 130
rect 919 1106 977 1118
rect 919 130 931 1106
rect 965 130 977 1106
rect 919 118 977 130
rect 1077 1106 1135 1118
rect 1077 130 1089 1106
rect 1123 130 1135 1106
rect 1077 118 1135 130
rect 1235 1106 1293 1118
rect 1235 130 1247 1106
rect 1281 130 1293 1106
rect 1235 118 1293 130
rect 1393 1106 1451 1118
rect 1393 130 1405 1106
rect 1439 130 1451 1106
rect 1393 118 1451 130
rect 1551 1106 1609 1118
rect 1551 130 1563 1106
rect 1597 130 1609 1106
rect 1551 118 1609 130
rect 1709 1106 1767 1118
rect 1709 130 1721 1106
rect 1755 130 1767 1106
rect 1709 118 1767 130
rect 1867 1106 1925 1118
rect 1867 130 1879 1106
rect 1913 130 1925 1106
rect 1867 118 1925 130
rect 2025 1106 2083 1118
rect 2025 130 2037 1106
rect 2071 130 2083 1106
rect 2025 118 2083 130
rect 2183 1106 2241 1118
rect 2183 130 2195 1106
rect 2229 130 2241 1106
rect 2183 118 2241 130
rect 2341 1106 2399 1118
rect 2341 130 2353 1106
rect 2387 130 2399 1106
rect 2341 118 2399 130
rect 2499 1106 2557 1118
rect 2499 130 2511 1106
rect 2545 130 2557 1106
rect 2499 118 2557 130
rect 2657 1106 2715 1118
rect 2657 130 2669 1106
rect 2703 130 2715 1106
rect 2657 118 2715 130
rect 2815 1106 2873 1118
rect 2815 130 2827 1106
rect 2861 130 2873 1106
rect 2815 118 2873 130
rect 2973 1106 3031 1118
rect 2973 130 2985 1106
rect 3019 130 3031 1106
rect 2973 118 3031 130
rect 3131 1106 3189 1118
rect 3131 130 3143 1106
rect 3177 130 3189 1106
rect 3131 118 3189 130
rect 3289 1106 3347 1118
rect 3289 130 3301 1106
rect 3335 130 3347 1106
rect 3289 118 3347 130
rect 3447 1106 3505 1118
rect 3447 130 3459 1106
rect 3493 130 3505 1106
rect 3447 118 3505 130
rect 3605 1106 3663 1118
rect 3605 130 3617 1106
rect 3651 130 3663 1106
rect 3605 118 3663 130
rect 3763 1106 3821 1118
rect 3763 130 3775 1106
rect 3809 130 3821 1106
rect 3763 118 3821 130
rect 3921 1106 3979 1118
rect 3921 130 3933 1106
rect 3967 130 3979 1106
rect 3921 118 3979 130
rect 4079 1106 4137 1118
rect 4079 130 4091 1106
rect 4125 130 4137 1106
rect 4079 118 4137 130
rect 4237 1106 4295 1118
rect 4237 130 4249 1106
rect 4283 130 4295 1106
rect 4237 118 4295 130
rect 4395 1106 4453 1118
rect 4395 130 4407 1106
rect 4441 130 4453 1106
rect 4395 118 4453 130
rect 4553 1106 4611 1118
rect 4553 130 4565 1106
rect 4599 130 4611 1106
rect 4553 118 4611 130
rect 4711 1106 4769 1118
rect 4711 130 4723 1106
rect 4757 130 4769 1106
rect 4711 118 4769 130
rect 4869 1106 4927 1118
rect 4869 130 4881 1106
rect 4915 130 4927 1106
rect 4869 118 4927 130
rect -4927 -130 -4869 -118
rect -4927 -1106 -4915 -130
rect -4881 -1106 -4869 -130
rect -4927 -1118 -4869 -1106
rect -4769 -130 -4711 -118
rect -4769 -1106 -4757 -130
rect -4723 -1106 -4711 -130
rect -4769 -1118 -4711 -1106
rect -4611 -130 -4553 -118
rect -4611 -1106 -4599 -130
rect -4565 -1106 -4553 -130
rect -4611 -1118 -4553 -1106
rect -4453 -130 -4395 -118
rect -4453 -1106 -4441 -130
rect -4407 -1106 -4395 -130
rect -4453 -1118 -4395 -1106
rect -4295 -130 -4237 -118
rect -4295 -1106 -4283 -130
rect -4249 -1106 -4237 -130
rect -4295 -1118 -4237 -1106
rect -4137 -130 -4079 -118
rect -4137 -1106 -4125 -130
rect -4091 -1106 -4079 -130
rect -4137 -1118 -4079 -1106
rect -3979 -130 -3921 -118
rect -3979 -1106 -3967 -130
rect -3933 -1106 -3921 -130
rect -3979 -1118 -3921 -1106
rect -3821 -130 -3763 -118
rect -3821 -1106 -3809 -130
rect -3775 -1106 -3763 -130
rect -3821 -1118 -3763 -1106
rect -3663 -130 -3605 -118
rect -3663 -1106 -3651 -130
rect -3617 -1106 -3605 -130
rect -3663 -1118 -3605 -1106
rect -3505 -130 -3447 -118
rect -3505 -1106 -3493 -130
rect -3459 -1106 -3447 -130
rect -3505 -1118 -3447 -1106
rect -3347 -130 -3289 -118
rect -3347 -1106 -3335 -130
rect -3301 -1106 -3289 -130
rect -3347 -1118 -3289 -1106
rect -3189 -130 -3131 -118
rect -3189 -1106 -3177 -130
rect -3143 -1106 -3131 -130
rect -3189 -1118 -3131 -1106
rect -3031 -130 -2973 -118
rect -3031 -1106 -3019 -130
rect -2985 -1106 -2973 -130
rect -3031 -1118 -2973 -1106
rect -2873 -130 -2815 -118
rect -2873 -1106 -2861 -130
rect -2827 -1106 -2815 -130
rect -2873 -1118 -2815 -1106
rect -2715 -130 -2657 -118
rect -2715 -1106 -2703 -130
rect -2669 -1106 -2657 -130
rect -2715 -1118 -2657 -1106
rect -2557 -130 -2499 -118
rect -2557 -1106 -2545 -130
rect -2511 -1106 -2499 -130
rect -2557 -1118 -2499 -1106
rect -2399 -130 -2341 -118
rect -2399 -1106 -2387 -130
rect -2353 -1106 -2341 -130
rect -2399 -1118 -2341 -1106
rect -2241 -130 -2183 -118
rect -2241 -1106 -2229 -130
rect -2195 -1106 -2183 -130
rect -2241 -1118 -2183 -1106
rect -2083 -130 -2025 -118
rect -2083 -1106 -2071 -130
rect -2037 -1106 -2025 -130
rect -2083 -1118 -2025 -1106
rect -1925 -130 -1867 -118
rect -1925 -1106 -1913 -130
rect -1879 -1106 -1867 -130
rect -1925 -1118 -1867 -1106
rect -1767 -130 -1709 -118
rect -1767 -1106 -1755 -130
rect -1721 -1106 -1709 -130
rect -1767 -1118 -1709 -1106
rect -1609 -130 -1551 -118
rect -1609 -1106 -1597 -130
rect -1563 -1106 -1551 -130
rect -1609 -1118 -1551 -1106
rect -1451 -130 -1393 -118
rect -1451 -1106 -1439 -130
rect -1405 -1106 -1393 -130
rect -1451 -1118 -1393 -1106
rect -1293 -130 -1235 -118
rect -1293 -1106 -1281 -130
rect -1247 -1106 -1235 -130
rect -1293 -1118 -1235 -1106
rect -1135 -130 -1077 -118
rect -1135 -1106 -1123 -130
rect -1089 -1106 -1077 -130
rect -1135 -1118 -1077 -1106
rect -977 -130 -919 -118
rect -977 -1106 -965 -130
rect -931 -1106 -919 -130
rect -977 -1118 -919 -1106
rect -819 -130 -761 -118
rect -819 -1106 -807 -130
rect -773 -1106 -761 -130
rect -819 -1118 -761 -1106
rect -661 -130 -603 -118
rect -661 -1106 -649 -130
rect -615 -1106 -603 -130
rect -661 -1118 -603 -1106
rect -503 -130 -445 -118
rect -503 -1106 -491 -130
rect -457 -1106 -445 -130
rect -503 -1118 -445 -1106
rect -345 -130 -287 -118
rect -345 -1106 -333 -130
rect -299 -1106 -287 -130
rect -345 -1118 -287 -1106
rect -187 -130 -129 -118
rect -187 -1106 -175 -130
rect -141 -1106 -129 -130
rect -187 -1118 -129 -1106
rect -29 -130 29 -118
rect -29 -1106 -17 -130
rect 17 -1106 29 -130
rect -29 -1118 29 -1106
rect 129 -130 187 -118
rect 129 -1106 141 -130
rect 175 -1106 187 -130
rect 129 -1118 187 -1106
rect 287 -130 345 -118
rect 287 -1106 299 -130
rect 333 -1106 345 -130
rect 287 -1118 345 -1106
rect 445 -130 503 -118
rect 445 -1106 457 -130
rect 491 -1106 503 -130
rect 445 -1118 503 -1106
rect 603 -130 661 -118
rect 603 -1106 615 -130
rect 649 -1106 661 -130
rect 603 -1118 661 -1106
rect 761 -130 819 -118
rect 761 -1106 773 -130
rect 807 -1106 819 -130
rect 761 -1118 819 -1106
rect 919 -130 977 -118
rect 919 -1106 931 -130
rect 965 -1106 977 -130
rect 919 -1118 977 -1106
rect 1077 -130 1135 -118
rect 1077 -1106 1089 -130
rect 1123 -1106 1135 -130
rect 1077 -1118 1135 -1106
rect 1235 -130 1293 -118
rect 1235 -1106 1247 -130
rect 1281 -1106 1293 -130
rect 1235 -1118 1293 -1106
rect 1393 -130 1451 -118
rect 1393 -1106 1405 -130
rect 1439 -1106 1451 -130
rect 1393 -1118 1451 -1106
rect 1551 -130 1609 -118
rect 1551 -1106 1563 -130
rect 1597 -1106 1609 -130
rect 1551 -1118 1609 -1106
rect 1709 -130 1767 -118
rect 1709 -1106 1721 -130
rect 1755 -1106 1767 -130
rect 1709 -1118 1767 -1106
rect 1867 -130 1925 -118
rect 1867 -1106 1879 -130
rect 1913 -1106 1925 -130
rect 1867 -1118 1925 -1106
rect 2025 -130 2083 -118
rect 2025 -1106 2037 -130
rect 2071 -1106 2083 -130
rect 2025 -1118 2083 -1106
rect 2183 -130 2241 -118
rect 2183 -1106 2195 -130
rect 2229 -1106 2241 -130
rect 2183 -1118 2241 -1106
rect 2341 -130 2399 -118
rect 2341 -1106 2353 -130
rect 2387 -1106 2399 -130
rect 2341 -1118 2399 -1106
rect 2499 -130 2557 -118
rect 2499 -1106 2511 -130
rect 2545 -1106 2557 -130
rect 2499 -1118 2557 -1106
rect 2657 -130 2715 -118
rect 2657 -1106 2669 -130
rect 2703 -1106 2715 -130
rect 2657 -1118 2715 -1106
rect 2815 -130 2873 -118
rect 2815 -1106 2827 -130
rect 2861 -1106 2873 -130
rect 2815 -1118 2873 -1106
rect 2973 -130 3031 -118
rect 2973 -1106 2985 -130
rect 3019 -1106 3031 -130
rect 2973 -1118 3031 -1106
rect 3131 -130 3189 -118
rect 3131 -1106 3143 -130
rect 3177 -1106 3189 -130
rect 3131 -1118 3189 -1106
rect 3289 -130 3347 -118
rect 3289 -1106 3301 -130
rect 3335 -1106 3347 -130
rect 3289 -1118 3347 -1106
rect 3447 -130 3505 -118
rect 3447 -1106 3459 -130
rect 3493 -1106 3505 -130
rect 3447 -1118 3505 -1106
rect 3605 -130 3663 -118
rect 3605 -1106 3617 -130
rect 3651 -1106 3663 -130
rect 3605 -1118 3663 -1106
rect 3763 -130 3821 -118
rect 3763 -1106 3775 -130
rect 3809 -1106 3821 -130
rect 3763 -1118 3821 -1106
rect 3921 -130 3979 -118
rect 3921 -1106 3933 -130
rect 3967 -1106 3979 -130
rect 3921 -1118 3979 -1106
rect 4079 -130 4137 -118
rect 4079 -1106 4091 -130
rect 4125 -1106 4137 -130
rect 4079 -1118 4137 -1106
rect 4237 -130 4295 -118
rect 4237 -1106 4249 -130
rect 4283 -1106 4295 -130
rect 4237 -1118 4295 -1106
rect 4395 -130 4453 -118
rect 4395 -1106 4407 -130
rect 4441 -1106 4453 -130
rect 4395 -1118 4453 -1106
rect 4553 -130 4611 -118
rect 4553 -1106 4565 -130
rect 4599 -1106 4611 -130
rect 4553 -1118 4611 -1106
rect 4711 -130 4769 -118
rect 4711 -1106 4723 -130
rect 4757 -1106 4769 -130
rect 4711 -1118 4769 -1106
rect 4869 -130 4927 -118
rect 4869 -1106 4881 -130
rect 4915 -1106 4927 -130
rect 4869 -1118 4927 -1106
rect -4927 -1366 -4869 -1354
rect -4927 -2342 -4915 -1366
rect -4881 -2342 -4869 -1366
rect -4927 -2354 -4869 -2342
rect -4769 -1366 -4711 -1354
rect -4769 -2342 -4757 -1366
rect -4723 -2342 -4711 -1366
rect -4769 -2354 -4711 -2342
rect -4611 -1366 -4553 -1354
rect -4611 -2342 -4599 -1366
rect -4565 -2342 -4553 -1366
rect -4611 -2354 -4553 -2342
rect -4453 -1366 -4395 -1354
rect -4453 -2342 -4441 -1366
rect -4407 -2342 -4395 -1366
rect -4453 -2354 -4395 -2342
rect -4295 -1366 -4237 -1354
rect -4295 -2342 -4283 -1366
rect -4249 -2342 -4237 -1366
rect -4295 -2354 -4237 -2342
rect -4137 -1366 -4079 -1354
rect -4137 -2342 -4125 -1366
rect -4091 -2342 -4079 -1366
rect -4137 -2354 -4079 -2342
rect -3979 -1366 -3921 -1354
rect -3979 -2342 -3967 -1366
rect -3933 -2342 -3921 -1366
rect -3979 -2354 -3921 -2342
rect -3821 -1366 -3763 -1354
rect -3821 -2342 -3809 -1366
rect -3775 -2342 -3763 -1366
rect -3821 -2354 -3763 -2342
rect -3663 -1366 -3605 -1354
rect -3663 -2342 -3651 -1366
rect -3617 -2342 -3605 -1366
rect -3663 -2354 -3605 -2342
rect -3505 -1366 -3447 -1354
rect -3505 -2342 -3493 -1366
rect -3459 -2342 -3447 -1366
rect -3505 -2354 -3447 -2342
rect -3347 -1366 -3289 -1354
rect -3347 -2342 -3335 -1366
rect -3301 -2342 -3289 -1366
rect -3347 -2354 -3289 -2342
rect -3189 -1366 -3131 -1354
rect -3189 -2342 -3177 -1366
rect -3143 -2342 -3131 -1366
rect -3189 -2354 -3131 -2342
rect -3031 -1366 -2973 -1354
rect -3031 -2342 -3019 -1366
rect -2985 -2342 -2973 -1366
rect -3031 -2354 -2973 -2342
rect -2873 -1366 -2815 -1354
rect -2873 -2342 -2861 -1366
rect -2827 -2342 -2815 -1366
rect -2873 -2354 -2815 -2342
rect -2715 -1366 -2657 -1354
rect -2715 -2342 -2703 -1366
rect -2669 -2342 -2657 -1366
rect -2715 -2354 -2657 -2342
rect -2557 -1366 -2499 -1354
rect -2557 -2342 -2545 -1366
rect -2511 -2342 -2499 -1366
rect -2557 -2354 -2499 -2342
rect -2399 -1366 -2341 -1354
rect -2399 -2342 -2387 -1366
rect -2353 -2342 -2341 -1366
rect -2399 -2354 -2341 -2342
rect -2241 -1366 -2183 -1354
rect -2241 -2342 -2229 -1366
rect -2195 -2342 -2183 -1366
rect -2241 -2354 -2183 -2342
rect -2083 -1366 -2025 -1354
rect -2083 -2342 -2071 -1366
rect -2037 -2342 -2025 -1366
rect -2083 -2354 -2025 -2342
rect -1925 -1366 -1867 -1354
rect -1925 -2342 -1913 -1366
rect -1879 -2342 -1867 -1366
rect -1925 -2354 -1867 -2342
rect -1767 -1366 -1709 -1354
rect -1767 -2342 -1755 -1366
rect -1721 -2342 -1709 -1366
rect -1767 -2354 -1709 -2342
rect -1609 -1366 -1551 -1354
rect -1609 -2342 -1597 -1366
rect -1563 -2342 -1551 -1366
rect -1609 -2354 -1551 -2342
rect -1451 -1366 -1393 -1354
rect -1451 -2342 -1439 -1366
rect -1405 -2342 -1393 -1366
rect -1451 -2354 -1393 -2342
rect -1293 -1366 -1235 -1354
rect -1293 -2342 -1281 -1366
rect -1247 -2342 -1235 -1366
rect -1293 -2354 -1235 -2342
rect -1135 -1366 -1077 -1354
rect -1135 -2342 -1123 -1366
rect -1089 -2342 -1077 -1366
rect -1135 -2354 -1077 -2342
rect -977 -1366 -919 -1354
rect -977 -2342 -965 -1366
rect -931 -2342 -919 -1366
rect -977 -2354 -919 -2342
rect -819 -1366 -761 -1354
rect -819 -2342 -807 -1366
rect -773 -2342 -761 -1366
rect -819 -2354 -761 -2342
rect -661 -1366 -603 -1354
rect -661 -2342 -649 -1366
rect -615 -2342 -603 -1366
rect -661 -2354 -603 -2342
rect -503 -1366 -445 -1354
rect -503 -2342 -491 -1366
rect -457 -2342 -445 -1366
rect -503 -2354 -445 -2342
rect -345 -1366 -287 -1354
rect -345 -2342 -333 -1366
rect -299 -2342 -287 -1366
rect -345 -2354 -287 -2342
rect -187 -1366 -129 -1354
rect -187 -2342 -175 -1366
rect -141 -2342 -129 -1366
rect -187 -2354 -129 -2342
rect -29 -1366 29 -1354
rect -29 -2342 -17 -1366
rect 17 -2342 29 -1366
rect -29 -2354 29 -2342
rect 129 -1366 187 -1354
rect 129 -2342 141 -1366
rect 175 -2342 187 -1366
rect 129 -2354 187 -2342
rect 287 -1366 345 -1354
rect 287 -2342 299 -1366
rect 333 -2342 345 -1366
rect 287 -2354 345 -2342
rect 445 -1366 503 -1354
rect 445 -2342 457 -1366
rect 491 -2342 503 -1366
rect 445 -2354 503 -2342
rect 603 -1366 661 -1354
rect 603 -2342 615 -1366
rect 649 -2342 661 -1366
rect 603 -2354 661 -2342
rect 761 -1366 819 -1354
rect 761 -2342 773 -1366
rect 807 -2342 819 -1366
rect 761 -2354 819 -2342
rect 919 -1366 977 -1354
rect 919 -2342 931 -1366
rect 965 -2342 977 -1366
rect 919 -2354 977 -2342
rect 1077 -1366 1135 -1354
rect 1077 -2342 1089 -1366
rect 1123 -2342 1135 -1366
rect 1077 -2354 1135 -2342
rect 1235 -1366 1293 -1354
rect 1235 -2342 1247 -1366
rect 1281 -2342 1293 -1366
rect 1235 -2354 1293 -2342
rect 1393 -1366 1451 -1354
rect 1393 -2342 1405 -1366
rect 1439 -2342 1451 -1366
rect 1393 -2354 1451 -2342
rect 1551 -1366 1609 -1354
rect 1551 -2342 1563 -1366
rect 1597 -2342 1609 -1366
rect 1551 -2354 1609 -2342
rect 1709 -1366 1767 -1354
rect 1709 -2342 1721 -1366
rect 1755 -2342 1767 -1366
rect 1709 -2354 1767 -2342
rect 1867 -1366 1925 -1354
rect 1867 -2342 1879 -1366
rect 1913 -2342 1925 -1366
rect 1867 -2354 1925 -2342
rect 2025 -1366 2083 -1354
rect 2025 -2342 2037 -1366
rect 2071 -2342 2083 -1366
rect 2025 -2354 2083 -2342
rect 2183 -1366 2241 -1354
rect 2183 -2342 2195 -1366
rect 2229 -2342 2241 -1366
rect 2183 -2354 2241 -2342
rect 2341 -1366 2399 -1354
rect 2341 -2342 2353 -1366
rect 2387 -2342 2399 -1366
rect 2341 -2354 2399 -2342
rect 2499 -1366 2557 -1354
rect 2499 -2342 2511 -1366
rect 2545 -2342 2557 -1366
rect 2499 -2354 2557 -2342
rect 2657 -1366 2715 -1354
rect 2657 -2342 2669 -1366
rect 2703 -2342 2715 -1366
rect 2657 -2354 2715 -2342
rect 2815 -1366 2873 -1354
rect 2815 -2342 2827 -1366
rect 2861 -2342 2873 -1366
rect 2815 -2354 2873 -2342
rect 2973 -1366 3031 -1354
rect 2973 -2342 2985 -1366
rect 3019 -2342 3031 -1366
rect 2973 -2354 3031 -2342
rect 3131 -1366 3189 -1354
rect 3131 -2342 3143 -1366
rect 3177 -2342 3189 -1366
rect 3131 -2354 3189 -2342
rect 3289 -1366 3347 -1354
rect 3289 -2342 3301 -1366
rect 3335 -2342 3347 -1366
rect 3289 -2354 3347 -2342
rect 3447 -1366 3505 -1354
rect 3447 -2342 3459 -1366
rect 3493 -2342 3505 -1366
rect 3447 -2354 3505 -2342
rect 3605 -1366 3663 -1354
rect 3605 -2342 3617 -1366
rect 3651 -2342 3663 -1366
rect 3605 -2354 3663 -2342
rect 3763 -1366 3821 -1354
rect 3763 -2342 3775 -1366
rect 3809 -2342 3821 -1366
rect 3763 -2354 3821 -2342
rect 3921 -1366 3979 -1354
rect 3921 -2342 3933 -1366
rect 3967 -2342 3979 -1366
rect 3921 -2354 3979 -2342
rect 4079 -1366 4137 -1354
rect 4079 -2342 4091 -1366
rect 4125 -2342 4137 -1366
rect 4079 -2354 4137 -2342
rect 4237 -1366 4295 -1354
rect 4237 -2342 4249 -1366
rect 4283 -2342 4295 -1366
rect 4237 -2354 4295 -2342
rect 4395 -1366 4453 -1354
rect 4395 -2342 4407 -1366
rect 4441 -2342 4453 -1366
rect 4395 -2354 4453 -2342
rect 4553 -1366 4611 -1354
rect 4553 -2342 4565 -1366
rect 4599 -2342 4611 -1366
rect 4553 -2354 4611 -2342
rect 4711 -1366 4769 -1354
rect 4711 -2342 4723 -1366
rect 4757 -2342 4769 -1366
rect 4711 -2354 4769 -2342
rect 4869 -1366 4927 -1354
rect 4869 -2342 4881 -1366
rect 4915 -2342 4927 -1366
rect 4869 -2354 4927 -2342
<< mvpdiffc >>
rect -4915 1366 -4881 2342
rect -4757 1366 -4723 2342
rect -4599 1366 -4565 2342
rect -4441 1366 -4407 2342
rect -4283 1366 -4249 2342
rect -4125 1366 -4091 2342
rect -3967 1366 -3933 2342
rect -3809 1366 -3775 2342
rect -3651 1366 -3617 2342
rect -3493 1366 -3459 2342
rect -3335 1366 -3301 2342
rect -3177 1366 -3143 2342
rect -3019 1366 -2985 2342
rect -2861 1366 -2827 2342
rect -2703 1366 -2669 2342
rect -2545 1366 -2511 2342
rect -2387 1366 -2353 2342
rect -2229 1366 -2195 2342
rect -2071 1366 -2037 2342
rect -1913 1366 -1879 2342
rect -1755 1366 -1721 2342
rect -1597 1366 -1563 2342
rect -1439 1366 -1405 2342
rect -1281 1366 -1247 2342
rect -1123 1366 -1089 2342
rect -965 1366 -931 2342
rect -807 1366 -773 2342
rect -649 1366 -615 2342
rect -491 1366 -457 2342
rect -333 1366 -299 2342
rect -175 1366 -141 2342
rect -17 1366 17 2342
rect 141 1366 175 2342
rect 299 1366 333 2342
rect 457 1366 491 2342
rect 615 1366 649 2342
rect 773 1366 807 2342
rect 931 1366 965 2342
rect 1089 1366 1123 2342
rect 1247 1366 1281 2342
rect 1405 1366 1439 2342
rect 1563 1366 1597 2342
rect 1721 1366 1755 2342
rect 1879 1366 1913 2342
rect 2037 1366 2071 2342
rect 2195 1366 2229 2342
rect 2353 1366 2387 2342
rect 2511 1366 2545 2342
rect 2669 1366 2703 2342
rect 2827 1366 2861 2342
rect 2985 1366 3019 2342
rect 3143 1366 3177 2342
rect 3301 1366 3335 2342
rect 3459 1366 3493 2342
rect 3617 1366 3651 2342
rect 3775 1366 3809 2342
rect 3933 1366 3967 2342
rect 4091 1366 4125 2342
rect 4249 1366 4283 2342
rect 4407 1366 4441 2342
rect 4565 1366 4599 2342
rect 4723 1366 4757 2342
rect 4881 1366 4915 2342
rect -4915 130 -4881 1106
rect -4757 130 -4723 1106
rect -4599 130 -4565 1106
rect -4441 130 -4407 1106
rect -4283 130 -4249 1106
rect -4125 130 -4091 1106
rect -3967 130 -3933 1106
rect -3809 130 -3775 1106
rect -3651 130 -3617 1106
rect -3493 130 -3459 1106
rect -3335 130 -3301 1106
rect -3177 130 -3143 1106
rect -3019 130 -2985 1106
rect -2861 130 -2827 1106
rect -2703 130 -2669 1106
rect -2545 130 -2511 1106
rect -2387 130 -2353 1106
rect -2229 130 -2195 1106
rect -2071 130 -2037 1106
rect -1913 130 -1879 1106
rect -1755 130 -1721 1106
rect -1597 130 -1563 1106
rect -1439 130 -1405 1106
rect -1281 130 -1247 1106
rect -1123 130 -1089 1106
rect -965 130 -931 1106
rect -807 130 -773 1106
rect -649 130 -615 1106
rect -491 130 -457 1106
rect -333 130 -299 1106
rect -175 130 -141 1106
rect -17 130 17 1106
rect 141 130 175 1106
rect 299 130 333 1106
rect 457 130 491 1106
rect 615 130 649 1106
rect 773 130 807 1106
rect 931 130 965 1106
rect 1089 130 1123 1106
rect 1247 130 1281 1106
rect 1405 130 1439 1106
rect 1563 130 1597 1106
rect 1721 130 1755 1106
rect 1879 130 1913 1106
rect 2037 130 2071 1106
rect 2195 130 2229 1106
rect 2353 130 2387 1106
rect 2511 130 2545 1106
rect 2669 130 2703 1106
rect 2827 130 2861 1106
rect 2985 130 3019 1106
rect 3143 130 3177 1106
rect 3301 130 3335 1106
rect 3459 130 3493 1106
rect 3617 130 3651 1106
rect 3775 130 3809 1106
rect 3933 130 3967 1106
rect 4091 130 4125 1106
rect 4249 130 4283 1106
rect 4407 130 4441 1106
rect 4565 130 4599 1106
rect 4723 130 4757 1106
rect 4881 130 4915 1106
rect -4915 -1106 -4881 -130
rect -4757 -1106 -4723 -130
rect -4599 -1106 -4565 -130
rect -4441 -1106 -4407 -130
rect -4283 -1106 -4249 -130
rect -4125 -1106 -4091 -130
rect -3967 -1106 -3933 -130
rect -3809 -1106 -3775 -130
rect -3651 -1106 -3617 -130
rect -3493 -1106 -3459 -130
rect -3335 -1106 -3301 -130
rect -3177 -1106 -3143 -130
rect -3019 -1106 -2985 -130
rect -2861 -1106 -2827 -130
rect -2703 -1106 -2669 -130
rect -2545 -1106 -2511 -130
rect -2387 -1106 -2353 -130
rect -2229 -1106 -2195 -130
rect -2071 -1106 -2037 -130
rect -1913 -1106 -1879 -130
rect -1755 -1106 -1721 -130
rect -1597 -1106 -1563 -130
rect -1439 -1106 -1405 -130
rect -1281 -1106 -1247 -130
rect -1123 -1106 -1089 -130
rect -965 -1106 -931 -130
rect -807 -1106 -773 -130
rect -649 -1106 -615 -130
rect -491 -1106 -457 -130
rect -333 -1106 -299 -130
rect -175 -1106 -141 -130
rect -17 -1106 17 -130
rect 141 -1106 175 -130
rect 299 -1106 333 -130
rect 457 -1106 491 -130
rect 615 -1106 649 -130
rect 773 -1106 807 -130
rect 931 -1106 965 -130
rect 1089 -1106 1123 -130
rect 1247 -1106 1281 -130
rect 1405 -1106 1439 -130
rect 1563 -1106 1597 -130
rect 1721 -1106 1755 -130
rect 1879 -1106 1913 -130
rect 2037 -1106 2071 -130
rect 2195 -1106 2229 -130
rect 2353 -1106 2387 -130
rect 2511 -1106 2545 -130
rect 2669 -1106 2703 -130
rect 2827 -1106 2861 -130
rect 2985 -1106 3019 -130
rect 3143 -1106 3177 -130
rect 3301 -1106 3335 -130
rect 3459 -1106 3493 -130
rect 3617 -1106 3651 -130
rect 3775 -1106 3809 -130
rect 3933 -1106 3967 -130
rect 4091 -1106 4125 -130
rect 4249 -1106 4283 -130
rect 4407 -1106 4441 -130
rect 4565 -1106 4599 -130
rect 4723 -1106 4757 -130
rect 4881 -1106 4915 -130
rect -4915 -2342 -4881 -1366
rect -4757 -2342 -4723 -1366
rect -4599 -2342 -4565 -1366
rect -4441 -2342 -4407 -1366
rect -4283 -2342 -4249 -1366
rect -4125 -2342 -4091 -1366
rect -3967 -2342 -3933 -1366
rect -3809 -2342 -3775 -1366
rect -3651 -2342 -3617 -1366
rect -3493 -2342 -3459 -1366
rect -3335 -2342 -3301 -1366
rect -3177 -2342 -3143 -1366
rect -3019 -2342 -2985 -1366
rect -2861 -2342 -2827 -1366
rect -2703 -2342 -2669 -1366
rect -2545 -2342 -2511 -1366
rect -2387 -2342 -2353 -1366
rect -2229 -2342 -2195 -1366
rect -2071 -2342 -2037 -1366
rect -1913 -2342 -1879 -1366
rect -1755 -2342 -1721 -1366
rect -1597 -2342 -1563 -1366
rect -1439 -2342 -1405 -1366
rect -1281 -2342 -1247 -1366
rect -1123 -2342 -1089 -1366
rect -965 -2342 -931 -1366
rect -807 -2342 -773 -1366
rect -649 -2342 -615 -1366
rect -491 -2342 -457 -1366
rect -333 -2342 -299 -1366
rect -175 -2342 -141 -1366
rect -17 -2342 17 -1366
rect 141 -2342 175 -1366
rect 299 -2342 333 -1366
rect 457 -2342 491 -1366
rect 615 -2342 649 -1366
rect 773 -2342 807 -1366
rect 931 -2342 965 -1366
rect 1089 -2342 1123 -1366
rect 1247 -2342 1281 -1366
rect 1405 -2342 1439 -1366
rect 1563 -2342 1597 -1366
rect 1721 -2342 1755 -1366
rect 1879 -2342 1913 -1366
rect 2037 -2342 2071 -1366
rect 2195 -2342 2229 -1366
rect 2353 -2342 2387 -1366
rect 2511 -2342 2545 -1366
rect 2669 -2342 2703 -1366
rect 2827 -2342 2861 -1366
rect 2985 -2342 3019 -1366
rect 3143 -2342 3177 -1366
rect 3301 -2342 3335 -1366
rect 3459 -2342 3493 -1366
rect 3617 -2342 3651 -1366
rect 3775 -2342 3809 -1366
rect 3933 -2342 3967 -1366
rect 4091 -2342 4125 -1366
rect 4249 -2342 4283 -1366
rect 4407 -2342 4441 -1366
rect 4565 -2342 4599 -1366
rect 4723 -2342 4757 -1366
rect 4881 -2342 4915 -1366
<< mvnsubdiff >>
rect -5061 2573 5061 2585
rect -5061 2539 -4953 2573
rect 4953 2539 5061 2573
rect -5061 2527 5061 2539
rect -5061 2477 -5003 2527
rect -5061 -2477 -5049 2477
rect -5015 -2477 -5003 2477
rect 5003 2477 5061 2527
rect -5061 -2527 -5003 -2477
rect 5003 -2477 5015 2477
rect 5049 -2477 5061 2477
rect 5003 -2527 5061 -2477
rect -5061 -2539 5061 -2527
rect -5061 -2573 -4953 -2539
rect 4953 -2573 5061 -2539
rect -5061 -2585 5061 -2573
<< mvnsubdiffcont >>
rect -4953 2539 4953 2573
rect -5049 -2477 -5015 2477
rect 5015 -2477 5049 2477
rect -4953 -2573 4953 -2539
<< poly >>
rect -4869 2435 -4769 2451
rect -4869 2401 -4853 2435
rect -4785 2401 -4769 2435
rect -4869 2354 -4769 2401
rect -4711 2435 -4611 2451
rect -4711 2401 -4695 2435
rect -4627 2401 -4611 2435
rect -4711 2354 -4611 2401
rect -4553 2435 -4453 2451
rect -4553 2401 -4537 2435
rect -4469 2401 -4453 2435
rect -4553 2354 -4453 2401
rect -4395 2435 -4295 2451
rect -4395 2401 -4379 2435
rect -4311 2401 -4295 2435
rect -4395 2354 -4295 2401
rect -4237 2435 -4137 2451
rect -4237 2401 -4221 2435
rect -4153 2401 -4137 2435
rect -4237 2354 -4137 2401
rect -4079 2435 -3979 2451
rect -4079 2401 -4063 2435
rect -3995 2401 -3979 2435
rect -4079 2354 -3979 2401
rect -3921 2435 -3821 2451
rect -3921 2401 -3905 2435
rect -3837 2401 -3821 2435
rect -3921 2354 -3821 2401
rect -3763 2435 -3663 2451
rect -3763 2401 -3747 2435
rect -3679 2401 -3663 2435
rect -3763 2354 -3663 2401
rect -3605 2435 -3505 2451
rect -3605 2401 -3589 2435
rect -3521 2401 -3505 2435
rect -3605 2354 -3505 2401
rect -3447 2435 -3347 2451
rect -3447 2401 -3431 2435
rect -3363 2401 -3347 2435
rect -3447 2354 -3347 2401
rect -3289 2435 -3189 2451
rect -3289 2401 -3273 2435
rect -3205 2401 -3189 2435
rect -3289 2354 -3189 2401
rect -3131 2435 -3031 2451
rect -3131 2401 -3115 2435
rect -3047 2401 -3031 2435
rect -3131 2354 -3031 2401
rect -2973 2435 -2873 2451
rect -2973 2401 -2957 2435
rect -2889 2401 -2873 2435
rect -2973 2354 -2873 2401
rect -2815 2435 -2715 2451
rect -2815 2401 -2799 2435
rect -2731 2401 -2715 2435
rect -2815 2354 -2715 2401
rect -2657 2435 -2557 2451
rect -2657 2401 -2641 2435
rect -2573 2401 -2557 2435
rect -2657 2354 -2557 2401
rect -2499 2435 -2399 2451
rect -2499 2401 -2483 2435
rect -2415 2401 -2399 2435
rect -2499 2354 -2399 2401
rect -2341 2435 -2241 2451
rect -2341 2401 -2325 2435
rect -2257 2401 -2241 2435
rect -2341 2354 -2241 2401
rect -2183 2435 -2083 2451
rect -2183 2401 -2167 2435
rect -2099 2401 -2083 2435
rect -2183 2354 -2083 2401
rect -2025 2435 -1925 2451
rect -2025 2401 -2009 2435
rect -1941 2401 -1925 2435
rect -2025 2354 -1925 2401
rect -1867 2435 -1767 2451
rect -1867 2401 -1851 2435
rect -1783 2401 -1767 2435
rect -1867 2354 -1767 2401
rect -1709 2435 -1609 2451
rect -1709 2401 -1693 2435
rect -1625 2401 -1609 2435
rect -1709 2354 -1609 2401
rect -1551 2435 -1451 2451
rect -1551 2401 -1535 2435
rect -1467 2401 -1451 2435
rect -1551 2354 -1451 2401
rect -1393 2435 -1293 2451
rect -1393 2401 -1377 2435
rect -1309 2401 -1293 2435
rect -1393 2354 -1293 2401
rect -1235 2435 -1135 2451
rect -1235 2401 -1219 2435
rect -1151 2401 -1135 2435
rect -1235 2354 -1135 2401
rect -1077 2435 -977 2451
rect -1077 2401 -1061 2435
rect -993 2401 -977 2435
rect -1077 2354 -977 2401
rect -919 2435 -819 2451
rect -919 2401 -903 2435
rect -835 2401 -819 2435
rect -919 2354 -819 2401
rect -761 2435 -661 2451
rect -761 2401 -745 2435
rect -677 2401 -661 2435
rect -761 2354 -661 2401
rect -603 2435 -503 2451
rect -603 2401 -587 2435
rect -519 2401 -503 2435
rect -603 2354 -503 2401
rect -445 2435 -345 2451
rect -445 2401 -429 2435
rect -361 2401 -345 2435
rect -445 2354 -345 2401
rect -287 2435 -187 2451
rect -287 2401 -271 2435
rect -203 2401 -187 2435
rect -287 2354 -187 2401
rect -129 2435 -29 2451
rect -129 2401 -113 2435
rect -45 2401 -29 2435
rect -129 2354 -29 2401
rect 29 2435 129 2451
rect 29 2401 45 2435
rect 113 2401 129 2435
rect 29 2354 129 2401
rect 187 2435 287 2451
rect 187 2401 203 2435
rect 271 2401 287 2435
rect 187 2354 287 2401
rect 345 2435 445 2451
rect 345 2401 361 2435
rect 429 2401 445 2435
rect 345 2354 445 2401
rect 503 2435 603 2451
rect 503 2401 519 2435
rect 587 2401 603 2435
rect 503 2354 603 2401
rect 661 2435 761 2451
rect 661 2401 677 2435
rect 745 2401 761 2435
rect 661 2354 761 2401
rect 819 2435 919 2451
rect 819 2401 835 2435
rect 903 2401 919 2435
rect 819 2354 919 2401
rect 977 2435 1077 2451
rect 977 2401 993 2435
rect 1061 2401 1077 2435
rect 977 2354 1077 2401
rect 1135 2435 1235 2451
rect 1135 2401 1151 2435
rect 1219 2401 1235 2435
rect 1135 2354 1235 2401
rect 1293 2435 1393 2451
rect 1293 2401 1309 2435
rect 1377 2401 1393 2435
rect 1293 2354 1393 2401
rect 1451 2435 1551 2451
rect 1451 2401 1467 2435
rect 1535 2401 1551 2435
rect 1451 2354 1551 2401
rect 1609 2435 1709 2451
rect 1609 2401 1625 2435
rect 1693 2401 1709 2435
rect 1609 2354 1709 2401
rect 1767 2435 1867 2451
rect 1767 2401 1783 2435
rect 1851 2401 1867 2435
rect 1767 2354 1867 2401
rect 1925 2435 2025 2451
rect 1925 2401 1941 2435
rect 2009 2401 2025 2435
rect 1925 2354 2025 2401
rect 2083 2435 2183 2451
rect 2083 2401 2099 2435
rect 2167 2401 2183 2435
rect 2083 2354 2183 2401
rect 2241 2435 2341 2451
rect 2241 2401 2257 2435
rect 2325 2401 2341 2435
rect 2241 2354 2341 2401
rect 2399 2435 2499 2451
rect 2399 2401 2415 2435
rect 2483 2401 2499 2435
rect 2399 2354 2499 2401
rect 2557 2435 2657 2451
rect 2557 2401 2573 2435
rect 2641 2401 2657 2435
rect 2557 2354 2657 2401
rect 2715 2435 2815 2451
rect 2715 2401 2731 2435
rect 2799 2401 2815 2435
rect 2715 2354 2815 2401
rect 2873 2435 2973 2451
rect 2873 2401 2889 2435
rect 2957 2401 2973 2435
rect 2873 2354 2973 2401
rect 3031 2435 3131 2451
rect 3031 2401 3047 2435
rect 3115 2401 3131 2435
rect 3031 2354 3131 2401
rect 3189 2435 3289 2451
rect 3189 2401 3205 2435
rect 3273 2401 3289 2435
rect 3189 2354 3289 2401
rect 3347 2435 3447 2451
rect 3347 2401 3363 2435
rect 3431 2401 3447 2435
rect 3347 2354 3447 2401
rect 3505 2435 3605 2451
rect 3505 2401 3521 2435
rect 3589 2401 3605 2435
rect 3505 2354 3605 2401
rect 3663 2435 3763 2451
rect 3663 2401 3679 2435
rect 3747 2401 3763 2435
rect 3663 2354 3763 2401
rect 3821 2435 3921 2451
rect 3821 2401 3837 2435
rect 3905 2401 3921 2435
rect 3821 2354 3921 2401
rect 3979 2435 4079 2451
rect 3979 2401 3995 2435
rect 4063 2401 4079 2435
rect 3979 2354 4079 2401
rect 4137 2435 4237 2451
rect 4137 2401 4153 2435
rect 4221 2401 4237 2435
rect 4137 2354 4237 2401
rect 4295 2435 4395 2451
rect 4295 2401 4311 2435
rect 4379 2401 4395 2435
rect 4295 2354 4395 2401
rect 4453 2435 4553 2451
rect 4453 2401 4469 2435
rect 4537 2401 4553 2435
rect 4453 2354 4553 2401
rect 4611 2435 4711 2451
rect 4611 2401 4627 2435
rect 4695 2401 4711 2435
rect 4611 2354 4711 2401
rect 4769 2435 4869 2451
rect 4769 2401 4785 2435
rect 4853 2401 4869 2435
rect 4769 2354 4869 2401
rect -4869 1307 -4769 1354
rect -4869 1273 -4853 1307
rect -4785 1273 -4769 1307
rect -4869 1257 -4769 1273
rect -4711 1307 -4611 1354
rect -4711 1273 -4695 1307
rect -4627 1273 -4611 1307
rect -4711 1257 -4611 1273
rect -4553 1307 -4453 1354
rect -4553 1273 -4537 1307
rect -4469 1273 -4453 1307
rect -4553 1257 -4453 1273
rect -4395 1307 -4295 1354
rect -4395 1273 -4379 1307
rect -4311 1273 -4295 1307
rect -4395 1257 -4295 1273
rect -4237 1307 -4137 1354
rect -4237 1273 -4221 1307
rect -4153 1273 -4137 1307
rect -4237 1257 -4137 1273
rect -4079 1307 -3979 1354
rect -4079 1273 -4063 1307
rect -3995 1273 -3979 1307
rect -4079 1257 -3979 1273
rect -3921 1307 -3821 1354
rect -3921 1273 -3905 1307
rect -3837 1273 -3821 1307
rect -3921 1257 -3821 1273
rect -3763 1307 -3663 1354
rect -3763 1273 -3747 1307
rect -3679 1273 -3663 1307
rect -3763 1257 -3663 1273
rect -3605 1307 -3505 1354
rect -3605 1273 -3589 1307
rect -3521 1273 -3505 1307
rect -3605 1257 -3505 1273
rect -3447 1307 -3347 1354
rect -3447 1273 -3431 1307
rect -3363 1273 -3347 1307
rect -3447 1257 -3347 1273
rect -3289 1307 -3189 1354
rect -3289 1273 -3273 1307
rect -3205 1273 -3189 1307
rect -3289 1257 -3189 1273
rect -3131 1307 -3031 1354
rect -3131 1273 -3115 1307
rect -3047 1273 -3031 1307
rect -3131 1257 -3031 1273
rect -2973 1307 -2873 1354
rect -2973 1273 -2957 1307
rect -2889 1273 -2873 1307
rect -2973 1257 -2873 1273
rect -2815 1307 -2715 1354
rect -2815 1273 -2799 1307
rect -2731 1273 -2715 1307
rect -2815 1257 -2715 1273
rect -2657 1307 -2557 1354
rect -2657 1273 -2641 1307
rect -2573 1273 -2557 1307
rect -2657 1257 -2557 1273
rect -2499 1307 -2399 1354
rect -2499 1273 -2483 1307
rect -2415 1273 -2399 1307
rect -2499 1257 -2399 1273
rect -2341 1307 -2241 1354
rect -2341 1273 -2325 1307
rect -2257 1273 -2241 1307
rect -2341 1257 -2241 1273
rect -2183 1307 -2083 1354
rect -2183 1273 -2167 1307
rect -2099 1273 -2083 1307
rect -2183 1257 -2083 1273
rect -2025 1307 -1925 1354
rect -2025 1273 -2009 1307
rect -1941 1273 -1925 1307
rect -2025 1257 -1925 1273
rect -1867 1307 -1767 1354
rect -1867 1273 -1851 1307
rect -1783 1273 -1767 1307
rect -1867 1257 -1767 1273
rect -1709 1307 -1609 1354
rect -1709 1273 -1693 1307
rect -1625 1273 -1609 1307
rect -1709 1257 -1609 1273
rect -1551 1307 -1451 1354
rect -1551 1273 -1535 1307
rect -1467 1273 -1451 1307
rect -1551 1257 -1451 1273
rect -1393 1307 -1293 1354
rect -1393 1273 -1377 1307
rect -1309 1273 -1293 1307
rect -1393 1257 -1293 1273
rect -1235 1307 -1135 1354
rect -1235 1273 -1219 1307
rect -1151 1273 -1135 1307
rect -1235 1257 -1135 1273
rect -1077 1307 -977 1354
rect -1077 1273 -1061 1307
rect -993 1273 -977 1307
rect -1077 1257 -977 1273
rect -919 1307 -819 1354
rect -919 1273 -903 1307
rect -835 1273 -819 1307
rect -919 1257 -819 1273
rect -761 1307 -661 1354
rect -761 1273 -745 1307
rect -677 1273 -661 1307
rect -761 1257 -661 1273
rect -603 1307 -503 1354
rect -603 1273 -587 1307
rect -519 1273 -503 1307
rect -603 1257 -503 1273
rect -445 1307 -345 1354
rect -445 1273 -429 1307
rect -361 1273 -345 1307
rect -445 1257 -345 1273
rect -287 1307 -187 1354
rect -287 1273 -271 1307
rect -203 1273 -187 1307
rect -287 1257 -187 1273
rect -129 1307 -29 1354
rect -129 1273 -113 1307
rect -45 1273 -29 1307
rect -129 1257 -29 1273
rect 29 1307 129 1354
rect 29 1273 45 1307
rect 113 1273 129 1307
rect 29 1257 129 1273
rect 187 1307 287 1354
rect 187 1273 203 1307
rect 271 1273 287 1307
rect 187 1257 287 1273
rect 345 1307 445 1354
rect 345 1273 361 1307
rect 429 1273 445 1307
rect 345 1257 445 1273
rect 503 1307 603 1354
rect 503 1273 519 1307
rect 587 1273 603 1307
rect 503 1257 603 1273
rect 661 1307 761 1354
rect 661 1273 677 1307
rect 745 1273 761 1307
rect 661 1257 761 1273
rect 819 1307 919 1354
rect 819 1273 835 1307
rect 903 1273 919 1307
rect 819 1257 919 1273
rect 977 1307 1077 1354
rect 977 1273 993 1307
rect 1061 1273 1077 1307
rect 977 1257 1077 1273
rect 1135 1307 1235 1354
rect 1135 1273 1151 1307
rect 1219 1273 1235 1307
rect 1135 1257 1235 1273
rect 1293 1307 1393 1354
rect 1293 1273 1309 1307
rect 1377 1273 1393 1307
rect 1293 1257 1393 1273
rect 1451 1307 1551 1354
rect 1451 1273 1467 1307
rect 1535 1273 1551 1307
rect 1451 1257 1551 1273
rect 1609 1307 1709 1354
rect 1609 1273 1625 1307
rect 1693 1273 1709 1307
rect 1609 1257 1709 1273
rect 1767 1307 1867 1354
rect 1767 1273 1783 1307
rect 1851 1273 1867 1307
rect 1767 1257 1867 1273
rect 1925 1307 2025 1354
rect 1925 1273 1941 1307
rect 2009 1273 2025 1307
rect 1925 1257 2025 1273
rect 2083 1307 2183 1354
rect 2083 1273 2099 1307
rect 2167 1273 2183 1307
rect 2083 1257 2183 1273
rect 2241 1307 2341 1354
rect 2241 1273 2257 1307
rect 2325 1273 2341 1307
rect 2241 1257 2341 1273
rect 2399 1307 2499 1354
rect 2399 1273 2415 1307
rect 2483 1273 2499 1307
rect 2399 1257 2499 1273
rect 2557 1307 2657 1354
rect 2557 1273 2573 1307
rect 2641 1273 2657 1307
rect 2557 1257 2657 1273
rect 2715 1307 2815 1354
rect 2715 1273 2731 1307
rect 2799 1273 2815 1307
rect 2715 1257 2815 1273
rect 2873 1307 2973 1354
rect 2873 1273 2889 1307
rect 2957 1273 2973 1307
rect 2873 1257 2973 1273
rect 3031 1307 3131 1354
rect 3031 1273 3047 1307
rect 3115 1273 3131 1307
rect 3031 1257 3131 1273
rect 3189 1307 3289 1354
rect 3189 1273 3205 1307
rect 3273 1273 3289 1307
rect 3189 1257 3289 1273
rect 3347 1307 3447 1354
rect 3347 1273 3363 1307
rect 3431 1273 3447 1307
rect 3347 1257 3447 1273
rect 3505 1307 3605 1354
rect 3505 1273 3521 1307
rect 3589 1273 3605 1307
rect 3505 1257 3605 1273
rect 3663 1307 3763 1354
rect 3663 1273 3679 1307
rect 3747 1273 3763 1307
rect 3663 1257 3763 1273
rect 3821 1307 3921 1354
rect 3821 1273 3837 1307
rect 3905 1273 3921 1307
rect 3821 1257 3921 1273
rect 3979 1307 4079 1354
rect 3979 1273 3995 1307
rect 4063 1273 4079 1307
rect 3979 1257 4079 1273
rect 4137 1307 4237 1354
rect 4137 1273 4153 1307
rect 4221 1273 4237 1307
rect 4137 1257 4237 1273
rect 4295 1307 4395 1354
rect 4295 1273 4311 1307
rect 4379 1273 4395 1307
rect 4295 1257 4395 1273
rect 4453 1307 4553 1354
rect 4453 1273 4469 1307
rect 4537 1273 4553 1307
rect 4453 1257 4553 1273
rect 4611 1307 4711 1354
rect 4611 1273 4627 1307
rect 4695 1273 4711 1307
rect 4611 1257 4711 1273
rect 4769 1307 4869 1354
rect 4769 1273 4785 1307
rect 4853 1273 4869 1307
rect 4769 1257 4869 1273
rect -4869 1199 -4769 1215
rect -4869 1165 -4853 1199
rect -4785 1165 -4769 1199
rect -4869 1118 -4769 1165
rect -4711 1199 -4611 1215
rect -4711 1165 -4695 1199
rect -4627 1165 -4611 1199
rect -4711 1118 -4611 1165
rect -4553 1199 -4453 1215
rect -4553 1165 -4537 1199
rect -4469 1165 -4453 1199
rect -4553 1118 -4453 1165
rect -4395 1199 -4295 1215
rect -4395 1165 -4379 1199
rect -4311 1165 -4295 1199
rect -4395 1118 -4295 1165
rect -4237 1199 -4137 1215
rect -4237 1165 -4221 1199
rect -4153 1165 -4137 1199
rect -4237 1118 -4137 1165
rect -4079 1199 -3979 1215
rect -4079 1165 -4063 1199
rect -3995 1165 -3979 1199
rect -4079 1118 -3979 1165
rect -3921 1199 -3821 1215
rect -3921 1165 -3905 1199
rect -3837 1165 -3821 1199
rect -3921 1118 -3821 1165
rect -3763 1199 -3663 1215
rect -3763 1165 -3747 1199
rect -3679 1165 -3663 1199
rect -3763 1118 -3663 1165
rect -3605 1199 -3505 1215
rect -3605 1165 -3589 1199
rect -3521 1165 -3505 1199
rect -3605 1118 -3505 1165
rect -3447 1199 -3347 1215
rect -3447 1165 -3431 1199
rect -3363 1165 -3347 1199
rect -3447 1118 -3347 1165
rect -3289 1199 -3189 1215
rect -3289 1165 -3273 1199
rect -3205 1165 -3189 1199
rect -3289 1118 -3189 1165
rect -3131 1199 -3031 1215
rect -3131 1165 -3115 1199
rect -3047 1165 -3031 1199
rect -3131 1118 -3031 1165
rect -2973 1199 -2873 1215
rect -2973 1165 -2957 1199
rect -2889 1165 -2873 1199
rect -2973 1118 -2873 1165
rect -2815 1199 -2715 1215
rect -2815 1165 -2799 1199
rect -2731 1165 -2715 1199
rect -2815 1118 -2715 1165
rect -2657 1199 -2557 1215
rect -2657 1165 -2641 1199
rect -2573 1165 -2557 1199
rect -2657 1118 -2557 1165
rect -2499 1199 -2399 1215
rect -2499 1165 -2483 1199
rect -2415 1165 -2399 1199
rect -2499 1118 -2399 1165
rect -2341 1199 -2241 1215
rect -2341 1165 -2325 1199
rect -2257 1165 -2241 1199
rect -2341 1118 -2241 1165
rect -2183 1199 -2083 1215
rect -2183 1165 -2167 1199
rect -2099 1165 -2083 1199
rect -2183 1118 -2083 1165
rect -2025 1199 -1925 1215
rect -2025 1165 -2009 1199
rect -1941 1165 -1925 1199
rect -2025 1118 -1925 1165
rect -1867 1199 -1767 1215
rect -1867 1165 -1851 1199
rect -1783 1165 -1767 1199
rect -1867 1118 -1767 1165
rect -1709 1199 -1609 1215
rect -1709 1165 -1693 1199
rect -1625 1165 -1609 1199
rect -1709 1118 -1609 1165
rect -1551 1199 -1451 1215
rect -1551 1165 -1535 1199
rect -1467 1165 -1451 1199
rect -1551 1118 -1451 1165
rect -1393 1199 -1293 1215
rect -1393 1165 -1377 1199
rect -1309 1165 -1293 1199
rect -1393 1118 -1293 1165
rect -1235 1199 -1135 1215
rect -1235 1165 -1219 1199
rect -1151 1165 -1135 1199
rect -1235 1118 -1135 1165
rect -1077 1199 -977 1215
rect -1077 1165 -1061 1199
rect -993 1165 -977 1199
rect -1077 1118 -977 1165
rect -919 1199 -819 1215
rect -919 1165 -903 1199
rect -835 1165 -819 1199
rect -919 1118 -819 1165
rect -761 1199 -661 1215
rect -761 1165 -745 1199
rect -677 1165 -661 1199
rect -761 1118 -661 1165
rect -603 1199 -503 1215
rect -603 1165 -587 1199
rect -519 1165 -503 1199
rect -603 1118 -503 1165
rect -445 1199 -345 1215
rect -445 1165 -429 1199
rect -361 1165 -345 1199
rect -445 1118 -345 1165
rect -287 1199 -187 1215
rect -287 1165 -271 1199
rect -203 1165 -187 1199
rect -287 1118 -187 1165
rect -129 1199 -29 1215
rect -129 1165 -113 1199
rect -45 1165 -29 1199
rect -129 1118 -29 1165
rect 29 1199 129 1215
rect 29 1165 45 1199
rect 113 1165 129 1199
rect 29 1118 129 1165
rect 187 1199 287 1215
rect 187 1165 203 1199
rect 271 1165 287 1199
rect 187 1118 287 1165
rect 345 1199 445 1215
rect 345 1165 361 1199
rect 429 1165 445 1199
rect 345 1118 445 1165
rect 503 1199 603 1215
rect 503 1165 519 1199
rect 587 1165 603 1199
rect 503 1118 603 1165
rect 661 1199 761 1215
rect 661 1165 677 1199
rect 745 1165 761 1199
rect 661 1118 761 1165
rect 819 1199 919 1215
rect 819 1165 835 1199
rect 903 1165 919 1199
rect 819 1118 919 1165
rect 977 1199 1077 1215
rect 977 1165 993 1199
rect 1061 1165 1077 1199
rect 977 1118 1077 1165
rect 1135 1199 1235 1215
rect 1135 1165 1151 1199
rect 1219 1165 1235 1199
rect 1135 1118 1235 1165
rect 1293 1199 1393 1215
rect 1293 1165 1309 1199
rect 1377 1165 1393 1199
rect 1293 1118 1393 1165
rect 1451 1199 1551 1215
rect 1451 1165 1467 1199
rect 1535 1165 1551 1199
rect 1451 1118 1551 1165
rect 1609 1199 1709 1215
rect 1609 1165 1625 1199
rect 1693 1165 1709 1199
rect 1609 1118 1709 1165
rect 1767 1199 1867 1215
rect 1767 1165 1783 1199
rect 1851 1165 1867 1199
rect 1767 1118 1867 1165
rect 1925 1199 2025 1215
rect 1925 1165 1941 1199
rect 2009 1165 2025 1199
rect 1925 1118 2025 1165
rect 2083 1199 2183 1215
rect 2083 1165 2099 1199
rect 2167 1165 2183 1199
rect 2083 1118 2183 1165
rect 2241 1199 2341 1215
rect 2241 1165 2257 1199
rect 2325 1165 2341 1199
rect 2241 1118 2341 1165
rect 2399 1199 2499 1215
rect 2399 1165 2415 1199
rect 2483 1165 2499 1199
rect 2399 1118 2499 1165
rect 2557 1199 2657 1215
rect 2557 1165 2573 1199
rect 2641 1165 2657 1199
rect 2557 1118 2657 1165
rect 2715 1199 2815 1215
rect 2715 1165 2731 1199
rect 2799 1165 2815 1199
rect 2715 1118 2815 1165
rect 2873 1199 2973 1215
rect 2873 1165 2889 1199
rect 2957 1165 2973 1199
rect 2873 1118 2973 1165
rect 3031 1199 3131 1215
rect 3031 1165 3047 1199
rect 3115 1165 3131 1199
rect 3031 1118 3131 1165
rect 3189 1199 3289 1215
rect 3189 1165 3205 1199
rect 3273 1165 3289 1199
rect 3189 1118 3289 1165
rect 3347 1199 3447 1215
rect 3347 1165 3363 1199
rect 3431 1165 3447 1199
rect 3347 1118 3447 1165
rect 3505 1199 3605 1215
rect 3505 1165 3521 1199
rect 3589 1165 3605 1199
rect 3505 1118 3605 1165
rect 3663 1199 3763 1215
rect 3663 1165 3679 1199
rect 3747 1165 3763 1199
rect 3663 1118 3763 1165
rect 3821 1199 3921 1215
rect 3821 1165 3837 1199
rect 3905 1165 3921 1199
rect 3821 1118 3921 1165
rect 3979 1199 4079 1215
rect 3979 1165 3995 1199
rect 4063 1165 4079 1199
rect 3979 1118 4079 1165
rect 4137 1199 4237 1215
rect 4137 1165 4153 1199
rect 4221 1165 4237 1199
rect 4137 1118 4237 1165
rect 4295 1199 4395 1215
rect 4295 1165 4311 1199
rect 4379 1165 4395 1199
rect 4295 1118 4395 1165
rect 4453 1199 4553 1215
rect 4453 1165 4469 1199
rect 4537 1165 4553 1199
rect 4453 1118 4553 1165
rect 4611 1199 4711 1215
rect 4611 1165 4627 1199
rect 4695 1165 4711 1199
rect 4611 1118 4711 1165
rect 4769 1199 4869 1215
rect 4769 1165 4785 1199
rect 4853 1165 4869 1199
rect 4769 1118 4869 1165
rect -4869 71 -4769 118
rect -4869 37 -4853 71
rect -4785 37 -4769 71
rect -4869 21 -4769 37
rect -4711 71 -4611 118
rect -4711 37 -4695 71
rect -4627 37 -4611 71
rect -4711 21 -4611 37
rect -4553 71 -4453 118
rect -4553 37 -4537 71
rect -4469 37 -4453 71
rect -4553 21 -4453 37
rect -4395 71 -4295 118
rect -4395 37 -4379 71
rect -4311 37 -4295 71
rect -4395 21 -4295 37
rect -4237 71 -4137 118
rect -4237 37 -4221 71
rect -4153 37 -4137 71
rect -4237 21 -4137 37
rect -4079 71 -3979 118
rect -4079 37 -4063 71
rect -3995 37 -3979 71
rect -4079 21 -3979 37
rect -3921 71 -3821 118
rect -3921 37 -3905 71
rect -3837 37 -3821 71
rect -3921 21 -3821 37
rect -3763 71 -3663 118
rect -3763 37 -3747 71
rect -3679 37 -3663 71
rect -3763 21 -3663 37
rect -3605 71 -3505 118
rect -3605 37 -3589 71
rect -3521 37 -3505 71
rect -3605 21 -3505 37
rect -3447 71 -3347 118
rect -3447 37 -3431 71
rect -3363 37 -3347 71
rect -3447 21 -3347 37
rect -3289 71 -3189 118
rect -3289 37 -3273 71
rect -3205 37 -3189 71
rect -3289 21 -3189 37
rect -3131 71 -3031 118
rect -3131 37 -3115 71
rect -3047 37 -3031 71
rect -3131 21 -3031 37
rect -2973 71 -2873 118
rect -2973 37 -2957 71
rect -2889 37 -2873 71
rect -2973 21 -2873 37
rect -2815 71 -2715 118
rect -2815 37 -2799 71
rect -2731 37 -2715 71
rect -2815 21 -2715 37
rect -2657 71 -2557 118
rect -2657 37 -2641 71
rect -2573 37 -2557 71
rect -2657 21 -2557 37
rect -2499 71 -2399 118
rect -2499 37 -2483 71
rect -2415 37 -2399 71
rect -2499 21 -2399 37
rect -2341 71 -2241 118
rect -2341 37 -2325 71
rect -2257 37 -2241 71
rect -2341 21 -2241 37
rect -2183 71 -2083 118
rect -2183 37 -2167 71
rect -2099 37 -2083 71
rect -2183 21 -2083 37
rect -2025 71 -1925 118
rect -2025 37 -2009 71
rect -1941 37 -1925 71
rect -2025 21 -1925 37
rect -1867 71 -1767 118
rect -1867 37 -1851 71
rect -1783 37 -1767 71
rect -1867 21 -1767 37
rect -1709 71 -1609 118
rect -1709 37 -1693 71
rect -1625 37 -1609 71
rect -1709 21 -1609 37
rect -1551 71 -1451 118
rect -1551 37 -1535 71
rect -1467 37 -1451 71
rect -1551 21 -1451 37
rect -1393 71 -1293 118
rect -1393 37 -1377 71
rect -1309 37 -1293 71
rect -1393 21 -1293 37
rect -1235 71 -1135 118
rect -1235 37 -1219 71
rect -1151 37 -1135 71
rect -1235 21 -1135 37
rect -1077 71 -977 118
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -1077 21 -977 37
rect -919 71 -819 118
rect -919 37 -903 71
rect -835 37 -819 71
rect -919 21 -819 37
rect -761 71 -661 118
rect -761 37 -745 71
rect -677 37 -661 71
rect -761 21 -661 37
rect -603 71 -503 118
rect -603 37 -587 71
rect -519 37 -503 71
rect -603 21 -503 37
rect -445 71 -345 118
rect -445 37 -429 71
rect -361 37 -345 71
rect -445 21 -345 37
rect -287 71 -187 118
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 118
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 118
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 118
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect 345 71 445 118
rect 345 37 361 71
rect 429 37 445 71
rect 345 21 445 37
rect 503 71 603 118
rect 503 37 519 71
rect 587 37 603 71
rect 503 21 603 37
rect 661 71 761 118
rect 661 37 677 71
rect 745 37 761 71
rect 661 21 761 37
rect 819 71 919 118
rect 819 37 835 71
rect 903 37 919 71
rect 819 21 919 37
rect 977 71 1077 118
rect 977 37 993 71
rect 1061 37 1077 71
rect 977 21 1077 37
rect 1135 71 1235 118
rect 1135 37 1151 71
rect 1219 37 1235 71
rect 1135 21 1235 37
rect 1293 71 1393 118
rect 1293 37 1309 71
rect 1377 37 1393 71
rect 1293 21 1393 37
rect 1451 71 1551 118
rect 1451 37 1467 71
rect 1535 37 1551 71
rect 1451 21 1551 37
rect 1609 71 1709 118
rect 1609 37 1625 71
rect 1693 37 1709 71
rect 1609 21 1709 37
rect 1767 71 1867 118
rect 1767 37 1783 71
rect 1851 37 1867 71
rect 1767 21 1867 37
rect 1925 71 2025 118
rect 1925 37 1941 71
rect 2009 37 2025 71
rect 1925 21 2025 37
rect 2083 71 2183 118
rect 2083 37 2099 71
rect 2167 37 2183 71
rect 2083 21 2183 37
rect 2241 71 2341 118
rect 2241 37 2257 71
rect 2325 37 2341 71
rect 2241 21 2341 37
rect 2399 71 2499 118
rect 2399 37 2415 71
rect 2483 37 2499 71
rect 2399 21 2499 37
rect 2557 71 2657 118
rect 2557 37 2573 71
rect 2641 37 2657 71
rect 2557 21 2657 37
rect 2715 71 2815 118
rect 2715 37 2731 71
rect 2799 37 2815 71
rect 2715 21 2815 37
rect 2873 71 2973 118
rect 2873 37 2889 71
rect 2957 37 2973 71
rect 2873 21 2973 37
rect 3031 71 3131 118
rect 3031 37 3047 71
rect 3115 37 3131 71
rect 3031 21 3131 37
rect 3189 71 3289 118
rect 3189 37 3205 71
rect 3273 37 3289 71
rect 3189 21 3289 37
rect 3347 71 3447 118
rect 3347 37 3363 71
rect 3431 37 3447 71
rect 3347 21 3447 37
rect 3505 71 3605 118
rect 3505 37 3521 71
rect 3589 37 3605 71
rect 3505 21 3605 37
rect 3663 71 3763 118
rect 3663 37 3679 71
rect 3747 37 3763 71
rect 3663 21 3763 37
rect 3821 71 3921 118
rect 3821 37 3837 71
rect 3905 37 3921 71
rect 3821 21 3921 37
rect 3979 71 4079 118
rect 3979 37 3995 71
rect 4063 37 4079 71
rect 3979 21 4079 37
rect 4137 71 4237 118
rect 4137 37 4153 71
rect 4221 37 4237 71
rect 4137 21 4237 37
rect 4295 71 4395 118
rect 4295 37 4311 71
rect 4379 37 4395 71
rect 4295 21 4395 37
rect 4453 71 4553 118
rect 4453 37 4469 71
rect 4537 37 4553 71
rect 4453 21 4553 37
rect 4611 71 4711 118
rect 4611 37 4627 71
rect 4695 37 4711 71
rect 4611 21 4711 37
rect 4769 71 4869 118
rect 4769 37 4785 71
rect 4853 37 4869 71
rect 4769 21 4869 37
rect -4869 -37 -4769 -21
rect -4869 -71 -4853 -37
rect -4785 -71 -4769 -37
rect -4869 -118 -4769 -71
rect -4711 -37 -4611 -21
rect -4711 -71 -4695 -37
rect -4627 -71 -4611 -37
rect -4711 -118 -4611 -71
rect -4553 -37 -4453 -21
rect -4553 -71 -4537 -37
rect -4469 -71 -4453 -37
rect -4553 -118 -4453 -71
rect -4395 -37 -4295 -21
rect -4395 -71 -4379 -37
rect -4311 -71 -4295 -37
rect -4395 -118 -4295 -71
rect -4237 -37 -4137 -21
rect -4237 -71 -4221 -37
rect -4153 -71 -4137 -37
rect -4237 -118 -4137 -71
rect -4079 -37 -3979 -21
rect -4079 -71 -4063 -37
rect -3995 -71 -3979 -37
rect -4079 -118 -3979 -71
rect -3921 -37 -3821 -21
rect -3921 -71 -3905 -37
rect -3837 -71 -3821 -37
rect -3921 -118 -3821 -71
rect -3763 -37 -3663 -21
rect -3763 -71 -3747 -37
rect -3679 -71 -3663 -37
rect -3763 -118 -3663 -71
rect -3605 -37 -3505 -21
rect -3605 -71 -3589 -37
rect -3521 -71 -3505 -37
rect -3605 -118 -3505 -71
rect -3447 -37 -3347 -21
rect -3447 -71 -3431 -37
rect -3363 -71 -3347 -37
rect -3447 -118 -3347 -71
rect -3289 -37 -3189 -21
rect -3289 -71 -3273 -37
rect -3205 -71 -3189 -37
rect -3289 -118 -3189 -71
rect -3131 -37 -3031 -21
rect -3131 -71 -3115 -37
rect -3047 -71 -3031 -37
rect -3131 -118 -3031 -71
rect -2973 -37 -2873 -21
rect -2973 -71 -2957 -37
rect -2889 -71 -2873 -37
rect -2973 -118 -2873 -71
rect -2815 -37 -2715 -21
rect -2815 -71 -2799 -37
rect -2731 -71 -2715 -37
rect -2815 -118 -2715 -71
rect -2657 -37 -2557 -21
rect -2657 -71 -2641 -37
rect -2573 -71 -2557 -37
rect -2657 -118 -2557 -71
rect -2499 -37 -2399 -21
rect -2499 -71 -2483 -37
rect -2415 -71 -2399 -37
rect -2499 -118 -2399 -71
rect -2341 -37 -2241 -21
rect -2341 -71 -2325 -37
rect -2257 -71 -2241 -37
rect -2341 -118 -2241 -71
rect -2183 -37 -2083 -21
rect -2183 -71 -2167 -37
rect -2099 -71 -2083 -37
rect -2183 -118 -2083 -71
rect -2025 -37 -1925 -21
rect -2025 -71 -2009 -37
rect -1941 -71 -1925 -37
rect -2025 -118 -1925 -71
rect -1867 -37 -1767 -21
rect -1867 -71 -1851 -37
rect -1783 -71 -1767 -37
rect -1867 -118 -1767 -71
rect -1709 -37 -1609 -21
rect -1709 -71 -1693 -37
rect -1625 -71 -1609 -37
rect -1709 -118 -1609 -71
rect -1551 -37 -1451 -21
rect -1551 -71 -1535 -37
rect -1467 -71 -1451 -37
rect -1551 -118 -1451 -71
rect -1393 -37 -1293 -21
rect -1393 -71 -1377 -37
rect -1309 -71 -1293 -37
rect -1393 -118 -1293 -71
rect -1235 -37 -1135 -21
rect -1235 -71 -1219 -37
rect -1151 -71 -1135 -37
rect -1235 -118 -1135 -71
rect -1077 -37 -977 -21
rect -1077 -71 -1061 -37
rect -993 -71 -977 -37
rect -1077 -118 -977 -71
rect -919 -37 -819 -21
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -919 -118 -819 -71
rect -761 -37 -661 -21
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -761 -118 -661 -71
rect -603 -37 -503 -21
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -603 -118 -503 -71
rect -445 -37 -345 -21
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -445 -118 -345 -71
rect -287 -37 -187 -21
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -287 -118 -187 -71
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -118 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -118 129 -71
rect 187 -37 287 -21
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 187 -118 287 -71
rect 345 -37 445 -21
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 345 -118 445 -71
rect 503 -37 603 -21
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 503 -118 603 -71
rect 661 -37 761 -21
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 661 -118 761 -71
rect 819 -37 919 -21
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 819 -118 919 -71
rect 977 -37 1077 -21
rect 977 -71 993 -37
rect 1061 -71 1077 -37
rect 977 -118 1077 -71
rect 1135 -37 1235 -21
rect 1135 -71 1151 -37
rect 1219 -71 1235 -37
rect 1135 -118 1235 -71
rect 1293 -37 1393 -21
rect 1293 -71 1309 -37
rect 1377 -71 1393 -37
rect 1293 -118 1393 -71
rect 1451 -37 1551 -21
rect 1451 -71 1467 -37
rect 1535 -71 1551 -37
rect 1451 -118 1551 -71
rect 1609 -37 1709 -21
rect 1609 -71 1625 -37
rect 1693 -71 1709 -37
rect 1609 -118 1709 -71
rect 1767 -37 1867 -21
rect 1767 -71 1783 -37
rect 1851 -71 1867 -37
rect 1767 -118 1867 -71
rect 1925 -37 2025 -21
rect 1925 -71 1941 -37
rect 2009 -71 2025 -37
rect 1925 -118 2025 -71
rect 2083 -37 2183 -21
rect 2083 -71 2099 -37
rect 2167 -71 2183 -37
rect 2083 -118 2183 -71
rect 2241 -37 2341 -21
rect 2241 -71 2257 -37
rect 2325 -71 2341 -37
rect 2241 -118 2341 -71
rect 2399 -37 2499 -21
rect 2399 -71 2415 -37
rect 2483 -71 2499 -37
rect 2399 -118 2499 -71
rect 2557 -37 2657 -21
rect 2557 -71 2573 -37
rect 2641 -71 2657 -37
rect 2557 -118 2657 -71
rect 2715 -37 2815 -21
rect 2715 -71 2731 -37
rect 2799 -71 2815 -37
rect 2715 -118 2815 -71
rect 2873 -37 2973 -21
rect 2873 -71 2889 -37
rect 2957 -71 2973 -37
rect 2873 -118 2973 -71
rect 3031 -37 3131 -21
rect 3031 -71 3047 -37
rect 3115 -71 3131 -37
rect 3031 -118 3131 -71
rect 3189 -37 3289 -21
rect 3189 -71 3205 -37
rect 3273 -71 3289 -37
rect 3189 -118 3289 -71
rect 3347 -37 3447 -21
rect 3347 -71 3363 -37
rect 3431 -71 3447 -37
rect 3347 -118 3447 -71
rect 3505 -37 3605 -21
rect 3505 -71 3521 -37
rect 3589 -71 3605 -37
rect 3505 -118 3605 -71
rect 3663 -37 3763 -21
rect 3663 -71 3679 -37
rect 3747 -71 3763 -37
rect 3663 -118 3763 -71
rect 3821 -37 3921 -21
rect 3821 -71 3837 -37
rect 3905 -71 3921 -37
rect 3821 -118 3921 -71
rect 3979 -37 4079 -21
rect 3979 -71 3995 -37
rect 4063 -71 4079 -37
rect 3979 -118 4079 -71
rect 4137 -37 4237 -21
rect 4137 -71 4153 -37
rect 4221 -71 4237 -37
rect 4137 -118 4237 -71
rect 4295 -37 4395 -21
rect 4295 -71 4311 -37
rect 4379 -71 4395 -37
rect 4295 -118 4395 -71
rect 4453 -37 4553 -21
rect 4453 -71 4469 -37
rect 4537 -71 4553 -37
rect 4453 -118 4553 -71
rect 4611 -37 4711 -21
rect 4611 -71 4627 -37
rect 4695 -71 4711 -37
rect 4611 -118 4711 -71
rect 4769 -37 4869 -21
rect 4769 -71 4785 -37
rect 4853 -71 4869 -37
rect 4769 -118 4869 -71
rect -4869 -1165 -4769 -1118
rect -4869 -1199 -4853 -1165
rect -4785 -1199 -4769 -1165
rect -4869 -1215 -4769 -1199
rect -4711 -1165 -4611 -1118
rect -4711 -1199 -4695 -1165
rect -4627 -1199 -4611 -1165
rect -4711 -1215 -4611 -1199
rect -4553 -1165 -4453 -1118
rect -4553 -1199 -4537 -1165
rect -4469 -1199 -4453 -1165
rect -4553 -1215 -4453 -1199
rect -4395 -1165 -4295 -1118
rect -4395 -1199 -4379 -1165
rect -4311 -1199 -4295 -1165
rect -4395 -1215 -4295 -1199
rect -4237 -1165 -4137 -1118
rect -4237 -1199 -4221 -1165
rect -4153 -1199 -4137 -1165
rect -4237 -1215 -4137 -1199
rect -4079 -1165 -3979 -1118
rect -4079 -1199 -4063 -1165
rect -3995 -1199 -3979 -1165
rect -4079 -1215 -3979 -1199
rect -3921 -1165 -3821 -1118
rect -3921 -1199 -3905 -1165
rect -3837 -1199 -3821 -1165
rect -3921 -1215 -3821 -1199
rect -3763 -1165 -3663 -1118
rect -3763 -1199 -3747 -1165
rect -3679 -1199 -3663 -1165
rect -3763 -1215 -3663 -1199
rect -3605 -1165 -3505 -1118
rect -3605 -1199 -3589 -1165
rect -3521 -1199 -3505 -1165
rect -3605 -1215 -3505 -1199
rect -3447 -1165 -3347 -1118
rect -3447 -1199 -3431 -1165
rect -3363 -1199 -3347 -1165
rect -3447 -1215 -3347 -1199
rect -3289 -1165 -3189 -1118
rect -3289 -1199 -3273 -1165
rect -3205 -1199 -3189 -1165
rect -3289 -1215 -3189 -1199
rect -3131 -1165 -3031 -1118
rect -3131 -1199 -3115 -1165
rect -3047 -1199 -3031 -1165
rect -3131 -1215 -3031 -1199
rect -2973 -1165 -2873 -1118
rect -2973 -1199 -2957 -1165
rect -2889 -1199 -2873 -1165
rect -2973 -1215 -2873 -1199
rect -2815 -1165 -2715 -1118
rect -2815 -1199 -2799 -1165
rect -2731 -1199 -2715 -1165
rect -2815 -1215 -2715 -1199
rect -2657 -1165 -2557 -1118
rect -2657 -1199 -2641 -1165
rect -2573 -1199 -2557 -1165
rect -2657 -1215 -2557 -1199
rect -2499 -1165 -2399 -1118
rect -2499 -1199 -2483 -1165
rect -2415 -1199 -2399 -1165
rect -2499 -1215 -2399 -1199
rect -2341 -1165 -2241 -1118
rect -2341 -1199 -2325 -1165
rect -2257 -1199 -2241 -1165
rect -2341 -1215 -2241 -1199
rect -2183 -1165 -2083 -1118
rect -2183 -1199 -2167 -1165
rect -2099 -1199 -2083 -1165
rect -2183 -1215 -2083 -1199
rect -2025 -1165 -1925 -1118
rect -2025 -1199 -2009 -1165
rect -1941 -1199 -1925 -1165
rect -2025 -1215 -1925 -1199
rect -1867 -1165 -1767 -1118
rect -1867 -1199 -1851 -1165
rect -1783 -1199 -1767 -1165
rect -1867 -1215 -1767 -1199
rect -1709 -1165 -1609 -1118
rect -1709 -1199 -1693 -1165
rect -1625 -1199 -1609 -1165
rect -1709 -1215 -1609 -1199
rect -1551 -1165 -1451 -1118
rect -1551 -1199 -1535 -1165
rect -1467 -1199 -1451 -1165
rect -1551 -1215 -1451 -1199
rect -1393 -1165 -1293 -1118
rect -1393 -1199 -1377 -1165
rect -1309 -1199 -1293 -1165
rect -1393 -1215 -1293 -1199
rect -1235 -1165 -1135 -1118
rect -1235 -1199 -1219 -1165
rect -1151 -1199 -1135 -1165
rect -1235 -1215 -1135 -1199
rect -1077 -1165 -977 -1118
rect -1077 -1199 -1061 -1165
rect -993 -1199 -977 -1165
rect -1077 -1215 -977 -1199
rect -919 -1165 -819 -1118
rect -919 -1199 -903 -1165
rect -835 -1199 -819 -1165
rect -919 -1215 -819 -1199
rect -761 -1165 -661 -1118
rect -761 -1199 -745 -1165
rect -677 -1199 -661 -1165
rect -761 -1215 -661 -1199
rect -603 -1165 -503 -1118
rect -603 -1199 -587 -1165
rect -519 -1199 -503 -1165
rect -603 -1215 -503 -1199
rect -445 -1165 -345 -1118
rect -445 -1199 -429 -1165
rect -361 -1199 -345 -1165
rect -445 -1215 -345 -1199
rect -287 -1165 -187 -1118
rect -287 -1199 -271 -1165
rect -203 -1199 -187 -1165
rect -287 -1215 -187 -1199
rect -129 -1165 -29 -1118
rect -129 -1199 -113 -1165
rect -45 -1199 -29 -1165
rect -129 -1215 -29 -1199
rect 29 -1165 129 -1118
rect 29 -1199 45 -1165
rect 113 -1199 129 -1165
rect 29 -1215 129 -1199
rect 187 -1165 287 -1118
rect 187 -1199 203 -1165
rect 271 -1199 287 -1165
rect 187 -1215 287 -1199
rect 345 -1165 445 -1118
rect 345 -1199 361 -1165
rect 429 -1199 445 -1165
rect 345 -1215 445 -1199
rect 503 -1165 603 -1118
rect 503 -1199 519 -1165
rect 587 -1199 603 -1165
rect 503 -1215 603 -1199
rect 661 -1165 761 -1118
rect 661 -1199 677 -1165
rect 745 -1199 761 -1165
rect 661 -1215 761 -1199
rect 819 -1165 919 -1118
rect 819 -1199 835 -1165
rect 903 -1199 919 -1165
rect 819 -1215 919 -1199
rect 977 -1165 1077 -1118
rect 977 -1199 993 -1165
rect 1061 -1199 1077 -1165
rect 977 -1215 1077 -1199
rect 1135 -1165 1235 -1118
rect 1135 -1199 1151 -1165
rect 1219 -1199 1235 -1165
rect 1135 -1215 1235 -1199
rect 1293 -1165 1393 -1118
rect 1293 -1199 1309 -1165
rect 1377 -1199 1393 -1165
rect 1293 -1215 1393 -1199
rect 1451 -1165 1551 -1118
rect 1451 -1199 1467 -1165
rect 1535 -1199 1551 -1165
rect 1451 -1215 1551 -1199
rect 1609 -1165 1709 -1118
rect 1609 -1199 1625 -1165
rect 1693 -1199 1709 -1165
rect 1609 -1215 1709 -1199
rect 1767 -1165 1867 -1118
rect 1767 -1199 1783 -1165
rect 1851 -1199 1867 -1165
rect 1767 -1215 1867 -1199
rect 1925 -1165 2025 -1118
rect 1925 -1199 1941 -1165
rect 2009 -1199 2025 -1165
rect 1925 -1215 2025 -1199
rect 2083 -1165 2183 -1118
rect 2083 -1199 2099 -1165
rect 2167 -1199 2183 -1165
rect 2083 -1215 2183 -1199
rect 2241 -1165 2341 -1118
rect 2241 -1199 2257 -1165
rect 2325 -1199 2341 -1165
rect 2241 -1215 2341 -1199
rect 2399 -1165 2499 -1118
rect 2399 -1199 2415 -1165
rect 2483 -1199 2499 -1165
rect 2399 -1215 2499 -1199
rect 2557 -1165 2657 -1118
rect 2557 -1199 2573 -1165
rect 2641 -1199 2657 -1165
rect 2557 -1215 2657 -1199
rect 2715 -1165 2815 -1118
rect 2715 -1199 2731 -1165
rect 2799 -1199 2815 -1165
rect 2715 -1215 2815 -1199
rect 2873 -1165 2973 -1118
rect 2873 -1199 2889 -1165
rect 2957 -1199 2973 -1165
rect 2873 -1215 2973 -1199
rect 3031 -1165 3131 -1118
rect 3031 -1199 3047 -1165
rect 3115 -1199 3131 -1165
rect 3031 -1215 3131 -1199
rect 3189 -1165 3289 -1118
rect 3189 -1199 3205 -1165
rect 3273 -1199 3289 -1165
rect 3189 -1215 3289 -1199
rect 3347 -1165 3447 -1118
rect 3347 -1199 3363 -1165
rect 3431 -1199 3447 -1165
rect 3347 -1215 3447 -1199
rect 3505 -1165 3605 -1118
rect 3505 -1199 3521 -1165
rect 3589 -1199 3605 -1165
rect 3505 -1215 3605 -1199
rect 3663 -1165 3763 -1118
rect 3663 -1199 3679 -1165
rect 3747 -1199 3763 -1165
rect 3663 -1215 3763 -1199
rect 3821 -1165 3921 -1118
rect 3821 -1199 3837 -1165
rect 3905 -1199 3921 -1165
rect 3821 -1215 3921 -1199
rect 3979 -1165 4079 -1118
rect 3979 -1199 3995 -1165
rect 4063 -1199 4079 -1165
rect 3979 -1215 4079 -1199
rect 4137 -1165 4237 -1118
rect 4137 -1199 4153 -1165
rect 4221 -1199 4237 -1165
rect 4137 -1215 4237 -1199
rect 4295 -1165 4395 -1118
rect 4295 -1199 4311 -1165
rect 4379 -1199 4395 -1165
rect 4295 -1215 4395 -1199
rect 4453 -1165 4553 -1118
rect 4453 -1199 4469 -1165
rect 4537 -1199 4553 -1165
rect 4453 -1215 4553 -1199
rect 4611 -1165 4711 -1118
rect 4611 -1199 4627 -1165
rect 4695 -1199 4711 -1165
rect 4611 -1215 4711 -1199
rect 4769 -1165 4869 -1118
rect 4769 -1199 4785 -1165
rect 4853 -1199 4869 -1165
rect 4769 -1215 4869 -1199
rect -4869 -1273 -4769 -1257
rect -4869 -1307 -4853 -1273
rect -4785 -1307 -4769 -1273
rect -4869 -1354 -4769 -1307
rect -4711 -1273 -4611 -1257
rect -4711 -1307 -4695 -1273
rect -4627 -1307 -4611 -1273
rect -4711 -1354 -4611 -1307
rect -4553 -1273 -4453 -1257
rect -4553 -1307 -4537 -1273
rect -4469 -1307 -4453 -1273
rect -4553 -1354 -4453 -1307
rect -4395 -1273 -4295 -1257
rect -4395 -1307 -4379 -1273
rect -4311 -1307 -4295 -1273
rect -4395 -1354 -4295 -1307
rect -4237 -1273 -4137 -1257
rect -4237 -1307 -4221 -1273
rect -4153 -1307 -4137 -1273
rect -4237 -1354 -4137 -1307
rect -4079 -1273 -3979 -1257
rect -4079 -1307 -4063 -1273
rect -3995 -1307 -3979 -1273
rect -4079 -1354 -3979 -1307
rect -3921 -1273 -3821 -1257
rect -3921 -1307 -3905 -1273
rect -3837 -1307 -3821 -1273
rect -3921 -1354 -3821 -1307
rect -3763 -1273 -3663 -1257
rect -3763 -1307 -3747 -1273
rect -3679 -1307 -3663 -1273
rect -3763 -1354 -3663 -1307
rect -3605 -1273 -3505 -1257
rect -3605 -1307 -3589 -1273
rect -3521 -1307 -3505 -1273
rect -3605 -1354 -3505 -1307
rect -3447 -1273 -3347 -1257
rect -3447 -1307 -3431 -1273
rect -3363 -1307 -3347 -1273
rect -3447 -1354 -3347 -1307
rect -3289 -1273 -3189 -1257
rect -3289 -1307 -3273 -1273
rect -3205 -1307 -3189 -1273
rect -3289 -1354 -3189 -1307
rect -3131 -1273 -3031 -1257
rect -3131 -1307 -3115 -1273
rect -3047 -1307 -3031 -1273
rect -3131 -1354 -3031 -1307
rect -2973 -1273 -2873 -1257
rect -2973 -1307 -2957 -1273
rect -2889 -1307 -2873 -1273
rect -2973 -1354 -2873 -1307
rect -2815 -1273 -2715 -1257
rect -2815 -1307 -2799 -1273
rect -2731 -1307 -2715 -1273
rect -2815 -1354 -2715 -1307
rect -2657 -1273 -2557 -1257
rect -2657 -1307 -2641 -1273
rect -2573 -1307 -2557 -1273
rect -2657 -1354 -2557 -1307
rect -2499 -1273 -2399 -1257
rect -2499 -1307 -2483 -1273
rect -2415 -1307 -2399 -1273
rect -2499 -1354 -2399 -1307
rect -2341 -1273 -2241 -1257
rect -2341 -1307 -2325 -1273
rect -2257 -1307 -2241 -1273
rect -2341 -1354 -2241 -1307
rect -2183 -1273 -2083 -1257
rect -2183 -1307 -2167 -1273
rect -2099 -1307 -2083 -1273
rect -2183 -1354 -2083 -1307
rect -2025 -1273 -1925 -1257
rect -2025 -1307 -2009 -1273
rect -1941 -1307 -1925 -1273
rect -2025 -1354 -1925 -1307
rect -1867 -1273 -1767 -1257
rect -1867 -1307 -1851 -1273
rect -1783 -1307 -1767 -1273
rect -1867 -1354 -1767 -1307
rect -1709 -1273 -1609 -1257
rect -1709 -1307 -1693 -1273
rect -1625 -1307 -1609 -1273
rect -1709 -1354 -1609 -1307
rect -1551 -1273 -1451 -1257
rect -1551 -1307 -1535 -1273
rect -1467 -1307 -1451 -1273
rect -1551 -1354 -1451 -1307
rect -1393 -1273 -1293 -1257
rect -1393 -1307 -1377 -1273
rect -1309 -1307 -1293 -1273
rect -1393 -1354 -1293 -1307
rect -1235 -1273 -1135 -1257
rect -1235 -1307 -1219 -1273
rect -1151 -1307 -1135 -1273
rect -1235 -1354 -1135 -1307
rect -1077 -1273 -977 -1257
rect -1077 -1307 -1061 -1273
rect -993 -1307 -977 -1273
rect -1077 -1354 -977 -1307
rect -919 -1273 -819 -1257
rect -919 -1307 -903 -1273
rect -835 -1307 -819 -1273
rect -919 -1354 -819 -1307
rect -761 -1273 -661 -1257
rect -761 -1307 -745 -1273
rect -677 -1307 -661 -1273
rect -761 -1354 -661 -1307
rect -603 -1273 -503 -1257
rect -603 -1307 -587 -1273
rect -519 -1307 -503 -1273
rect -603 -1354 -503 -1307
rect -445 -1273 -345 -1257
rect -445 -1307 -429 -1273
rect -361 -1307 -345 -1273
rect -445 -1354 -345 -1307
rect -287 -1273 -187 -1257
rect -287 -1307 -271 -1273
rect -203 -1307 -187 -1273
rect -287 -1354 -187 -1307
rect -129 -1273 -29 -1257
rect -129 -1307 -113 -1273
rect -45 -1307 -29 -1273
rect -129 -1354 -29 -1307
rect 29 -1273 129 -1257
rect 29 -1307 45 -1273
rect 113 -1307 129 -1273
rect 29 -1354 129 -1307
rect 187 -1273 287 -1257
rect 187 -1307 203 -1273
rect 271 -1307 287 -1273
rect 187 -1354 287 -1307
rect 345 -1273 445 -1257
rect 345 -1307 361 -1273
rect 429 -1307 445 -1273
rect 345 -1354 445 -1307
rect 503 -1273 603 -1257
rect 503 -1307 519 -1273
rect 587 -1307 603 -1273
rect 503 -1354 603 -1307
rect 661 -1273 761 -1257
rect 661 -1307 677 -1273
rect 745 -1307 761 -1273
rect 661 -1354 761 -1307
rect 819 -1273 919 -1257
rect 819 -1307 835 -1273
rect 903 -1307 919 -1273
rect 819 -1354 919 -1307
rect 977 -1273 1077 -1257
rect 977 -1307 993 -1273
rect 1061 -1307 1077 -1273
rect 977 -1354 1077 -1307
rect 1135 -1273 1235 -1257
rect 1135 -1307 1151 -1273
rect 1219 -1307 1235 -1273
rect 1135 -1354 1235 -1307
rect 1293 -1273 1393 -1257
rect 1293 -1307 1309 -1273
rect 1377 -1307 1393 -1273
rect 1293 -1354 1393 -1307
rect 1451 -1273 1551 -1257
rect 1451 -1307 1467 -1273
rect 1535 -1307 1551 -1273
rect 1451 -1354 1551 -1307
rect 1609 -1273 1709 -1257
rect 1609 -1307 1625 -1273
rect 1693 -1307 1709 -1273
rect 1609 -1354 1709 -1307
rect 1767 -1273 1867 -1257
rect 1767 -1307 1783 -1273
rect 1851 -1307 1867 -1273
rect 1767 -1354 1867 -1307
rect 1925 -1273 2025 -1257
rect 1925 -1307 1941 -1273
rect 2009 -1307 2025 -1273
rect 1925 -1354 2025 -1307
rect 2083 -1273 2183 -1257
rect 2083 -1307 2099 -1273
rect 2167 -1307 2183 -1273
rect 2083 -1354 2183 -1307
rect 2241 -1273 2341 -1257
rect 2241 -1307 2257 -1273
rect 2325 -1307 2341 -1273
rect 2241 -1354 2341 -1307
rect 2399 -1273 2499 -1257
rect 2399 -1307 2415 -1273
rect 2483 -1307 2499 -1273
rect 2399 -1354 2499 -1307
rect 2557 -1273 2657 -1257
rect 2557 -1307 2573 -1273
rect 2641 -1307 2657 -1273
rect 2557 -1354 2657 -1307
rect 2715 -1273 2815 -1257
rect 2715 -1307 2731 -1273
rect 2799 -1307 2815 -1273
rect 2715 -1354 2815 -1307
rect 2873 -1273 2973 -1257
rect 2873 -1307 2889 -1273
rect 2957 -1307 2973 -1273
rect 2873 -1354 2973 -1307
rect 3031 -1273 3131 -1257
rect 3031 -1307 3047 -1273
rect 3115 -1307 3131 -1273
rect 3031 -1354 3131 -1307
rect 3189 -1273 3289 -1257
rect 3189 -1307 3205 -1273
rect 3273 -1307 3289 -1273
rect 3189 -1354 3289 -1307
rect 3347 -1273 3447 -1257
rect 3347 -1307 3363 -1273
rect 3431 -1307 3447 -1273
rect 3347 -1354 3447 -1307
rect 3505 -1273 3605 -1257
rect 3505 -1307 3521 -1273
rect 3589 -1307 3605 -1273
rect 3505 -1354 3605 -1307
rect 3663 -1273 3763 -1257
rect 3663 -1307 3679 -1273
rect 3747 -1307 3763 -1273
rect 3663 -1354 3763 -1307
rect 3821 -1273 3921 -1257
rect 3821 -1307 3837 -1273
rect 3905 -1307 3921 -1273
rect 3821 -1354 3921 -1307
rect 3979 -1273 4079 -1257
rect 3979 -1307 3995 -1273
rect 4063 -1307 4079 -1273
rect 3979 -1354 4079 -1307
rect 4137 -1273 4237 -1257
rect 4137 -1307 4153 -1273
rect 4221 -1307 4237 -1273
rect 4137 -1354 4237 -1307
rect 4295 -1273 4395 -1257
rect 4295 -1307 4311 -1273
rect 4379 -1307 4395 -1273
rect 4295 -1354 4395 -1307
rect 4453 -1273 4553 -1257
rect 4453 -1307 4469 -1273
rect 4537 -1307 4553 -1273
rect 4453 -1354 4553 -1307
rect 4611 -1273 4711 -1257
rect 4611 -1307 4627 -1273
rect 4695 -1307 4711 -1273
rect 4611 -1354 4711 -1307
rect 4769 -1273 4869 -1257
rect 4769 -1307 4785 -1273
rect 4853 -1307 4869 -1273
rect 4769 -1354 4869 -1307
rect -4869 -2401 -4769 -2354
rect -4869 -2435 -4853 -2401
rect -4785 -2435 -4769 -2401
rect -4869 -2451 -4769 -2435
rect -4711 -2401 -4611 -2354
rect -4711 -2435 -4695 -2401
rect -4627 -2435 -4611 -2401
rect -4711 -2451 -4611 -2435
rect -4553 -2401 -4453 -2354
rect -4553 -2435 -4537 -2401
rect -4469 -2435 -4453 -2401
rect -4553 -2451 -4453 -2435
rect -4395 -2401 -4295 -2354
rect -4395 -2435 -4379 -2401
rect -4311 -2435 -4295 -2401
rect -4395 -2451 -4295 -2435
rect -4237 -2401 -4137 -2354
rect -4237 -2435 -4221 -2401
rect -4153 -2435 -4137 -2401
rect -4237 -2451 -4137 -2435
rect -4079 -2401 -3979 -2354
rect -4079 -2435 -4063 -2401
rect -3995 -2435 -3979 -2401
rect -4079 -2451 -3979 -2435
rect -3921 -2401 -3821 -2354
rect -3921 -2435 -3905 -2401
rect -3837 -2435 -3821 -2401
rect -3921 -2451 -3821 -2435
rect -3763 -2401 -3663 -2354
rect -3763 -2435 -3747 -2401
rect -3679 -2435 -3663 -2401
rect -3763 -2451 -3663 -2435
rect -3605 -2401 -3505 -2354
rect -3605 -2435 -3589 -2401
rect -3521 -2435 -3505 -2401
rect -3605 -2451 -3505 -2435
rect -3447 -2401 -3347 -2354
rect -3447 -2435 -3431 -2401
rect -3363 -2435 -3347 -2401
rect -3447 -2451 -3347 -2435
rect -3289 -2401 -3189 -2354
rect -3289 -2435 -3273 -2401
rect -3205 -2435 -3189 -2401
rect -3289 -2451 -3189 -2435
rect -3131 -2401 -3031 -2354
rect -3131 -2435 -3115 -2401
rect -3047 -2435 -3031 -2401
rect -3131 -2451 -3031 -2435
rect -2973 -2401 -2873 -2354
rect -2973 -2435 -2957 -2401
rect -2889 -2435 -2873 -2401
rect -2973 -2451 -2873 -2435
rect -2815 -2401 -2715 -2354
rect -2815 -2435 -2799 -2401
rect -2731 -2435 -2715 -2401
rect -2815 -2451 -2715 -2435
rect -2657 -2401 -2557 -2354
rect -2657 -2435 -2641 -2401
rect -2573 -2435 -2557 -2401
rect -2657 -2451 -2557 -2435
rect -2499 -2401 -2399 -2354
rect -2499 -2435 -2483 -2401
rect -2415 -2435 -2399 -2401
rect -2499 -2451 -2399 -2435
rect -2341 -2401 -2241 -2354
rect -2341 -2435 -2325 -2401
rect -2257 -2435 -2241 -2401
rect -2341 -2451 -2241 -2435
rect -2183 -2401 -2083 -2354
rect -2183 -2435 -2167 -2401
rect -2099 -2435 -2083 -2401
rect -2183 -2451 -2083 -2435
rect -2025 -2401 -1925 -2354
rect -2025 -2435 -2009 -2401
rect -1941 -2435 -1925 -2401
rect -2025 -2451 -1925 -2435
rect -1867 -2401 -1767 -2354
rect -1867 -2435 -1851 -2401
rect -1783 -2435 -1767 -2401
rect -1867 -2451 -1767 -2435
rect -1709 -2401 -1609 -2354
rect -1709 -2435 -1693 -2401
rect -1625 -2435 -1609 -2401
rect -1709 -2451 -1609 -2435
rect -1551 -2401 -1451 -2354
rect -1551 -2435 -1535 -2401
rect -1467 -2435 -1451 -2401
rect -1551 -2451 -1451 -2435
rect -1393 -2401 -1293 -2354
rect -1393 -2435 -1377 -2401
rect -1309 -2435 -1293 -2401
rect -1393 -2451 -1293 -2435
rect -1235 -2401 -1135 -2354
rect -1235 -2435 -1219 -2401
rect -1151 -2435 -1135 -2401
rect -1235 -2451 -1135 -2435
rect -1077 -2401 -977 -2354
rect -1077 -2435 -1061 -2401
rect -993 -2435 -977 -2401
rect -1077 -2451 -977 -2435
rect -919 -2401 -819 -2354
rect -919 -2435 -903 -2401
rect -835 -2435 -819 -2401
rect -919 -2451 -819 -2435
rect -761 -2401 -661 -2354
rect -761 -2435 -745 -2401
rect -677 -2435 -661 -2401
rect -761 -2451 -661 -2435
rect -603 -2401 -503 -2354
rect -603 -2435 -587 -2401
rect -519 -2435 -503 -2401
rect -603 -2451 -503 -2435
rect -445 -2401 -345 -2354
rect -445 -2435 -429 -2401
rect -361 -2435 -345 -2401
rect -445 -2451 -345 -2435
rect -287 -2401 -187 -2354
rect -287 -2435 -271 -2401
rect -203 -2435 -187 -2401
rect -287 -2451 -187 -2435
rect -129 -2401 -29 -2354
rect -129 -2435 -113 -2401
rect -45 -2435 -29 -2401
rect -129 -2451 -29 -2435
rect 29 -2401 129 -2354
rect 29 -2435 45 -2401
rect 113 -2435 129 -2401
rect 29 -2451 129 -2435
rect 187 -2401 287 -2354
rect 187 -2435 203 -2401
rect 271 -2435 287 -2401
rect 187 -2451 287 -2435
rect 345 -2401 445 -2354
rect 345 -2435 361 -2401
rect 429 -2435 445 -2401
rect 345 -2451 445 -2435
rect 503 -2401 603 -2354
rect 503 -2435 519 -2401
rect 587 -2435 603 -2401
rect 503 -2451 603 -2435
rect 661 -2401 761 -2354
rect 661 -2435 677 -2401
rect 745 -2435 761 -2401
rect 661 -2451 761 -2435
rect 819 -2401 919 -2354
rect 819 -2435 835 -2401
rect 903 -2435 919 -2401
rect 819 -2451 919 -2435
rect 977 -2401 1077 -2354
rect 977 -2435 993 -2401
rect 1061 -2435 1077 -2401
rect 977 -2451 1077 -2435
rect 1135 -2401 1235 -2354
rect 1135 -2435 1151 -2401
rect 1219 -2435 1235 -2401
rect 1135 -2451 1235 -2435
rect 1293 -2401 1393 -2354
rect 1293 -2435 1309 -2401
rect 1377 -2435 1393 -2401
rect 1293 -2451 1393 -2435
rect 1451 -2401 1551 -2354
rect 1451 -2435 1467 -2401
rect 1535 -2435 1551 -2401
rect 1451 -2451 1551 -2435
rect 1609 -2401 1709 -2354
rect 1609 -2435 1625 -2401
rect 1693 -2435 1709 -2401
rect 1609 -2451 1709 -2435
rect 1767 -2401 1867 -2354
rect 1767 -2435 1783 -2401
rect 1851 -2435 1867 -2401
rect 1767 -2451 1867 -2435
rect 1925 -2401 2025 -2354
rect 1925 -2435 1941 -2401
rect 2009 -2435 2025 -2401
rect 1925 -2451 2025 -2435
rect 2083 -2401 2183 -2354
rect 2083 -2435 2099 -2401
rect 2167 -2435 2183 -2401
rect 2083 -2451 2183 -2435
rect 2241 -2401 2341 -2354
rect 2241 -2435 2257 -2401
rect 2325 -2435 2341 -2401
rect 2241 -2451 2341 -2435
rect 2399 -2401 2499 -2354
rect 2399 -2435 2415 -2401
rect 2483 -2435 2499 -2401
rect 2399 -2451 2499 -2435
rect 2557 -2401 2657 -2354
rect 2557 -2435 2573 -2401
rect 2641 -2435 2657 -2401
rect 2557 -2451 2657 -2435
rect 2715 -2401 2815 -2354
rect 2715 -2435 2731 -2401
rect 2799 -2435 2815 -2401
rect 2715 -2451 2815 -2435
rect 2873 -2401 2973 -2354
rect 2873 -2435 2889 -2401
rect 2957 -2435 2973 -2401
rect 2873 -2451 2973 -2435
rect 3031 -2401 3131 -2354
rect 3031 -2435 3047 -2401
rect 3115 -2435 3131 -2401
rect 3031 -2451 3131 -2435
rect 3189 -2401 3289 -2354
rect 3189 -2435 3205 -2401
rect 3273 -2435 3289 -2401
rect 3189 -2451 3289 -2435
rect 3347 -2401 3447 -2354
rect 3347 -2435 3363 -2401
rect 3431 -2435 3447 -2401
rect 3347 -2451 3447 -2435
rect 3505 -2401 3605 -2354
rect 3505 -2435 3521 -2401
rect 3589 -2435 3605 -2401
rect 3505 -2451 3605 -2435
rect 3663 -2401 3763 -2354
rect 3663 -2435 3679 -2401
rect 3747 -2435 3763 -2401
rect 3663 -2451 3763 -2435
rect 3821 -2401 3921 -2354
rect 3821 -2435 3837 -2401
rect 3905 -2435 3921 -2401
rect 3821 -2451 3921 -2435
rect 3979 -2401 4079 -2354
rect 3979 -2435 3995 -2401
rect 4063 -2435 4079 -2401
rect 3979 -2451 4079 -2435
rect 4137 -2401 4237 -2354
rect 4137 -2435 4153 -2401
rect 4221 -2435 4237 -2401
rect 4137 -2451 4237 -2435
rect 4295 -2401 4395 -2354
rect 4295 -2435 4311 -2401
rect 4379 -2435 4395 -2401
rect 4295 -2451 4395 -2435
rect 4453 -2401 4553 -2354
rect 4453 -2435 4469 -2401
rect 4537 -2435 4553 -2401
rect 4453 -2451 4553 -2435
rect 4611 -2401 4711 -2354
rect 4611 -2435 4627 -2401
rect 4695 -2435 4711 -2401
rect 4611 -2451 4711 -2435
rect 4769 -2401 4869 -2354
rect 4769 -2435 4785 -2401
rect 4853 -2435 4869 -2401
rect 4769 -2451 4869 -2435
<< polycont >>
rect -4853 2401 -4785 2435
rect -4695 2401 -4627 2435
rect -4537 2401 -4469 2435
rect -4379 2401 -4311 2435
rect -4221 2401 -4153 2435
rect -4063 2401 -3995 2435
rect -3905 2401 -3837 2435
rect -3747 2401 -3679 2435
rect -3589 2401 -3521 2435
rect -3431 2401 -3363 2435
rect -3273 2401 -3205 2435
rect -3115 2401 -3047 2435
rect -2957 2401 -2889 2435
rect -2799 2401 -2731 2435
rect -2641 2401 -2573 2435
rect -2483 2401 -2415 2435
rect -2325 2401 -2257 2435
rect -2167 2401 -2099 2435
rect -2009 2401 -1941 2435
rect -1851 2401 -1783 2435
rect -1693 2401 -1625 2435
rect -1535 2401 -1467 2435
rect -1377 2401 -1309 2435
rect -1219 2401 -1151 2435
rect -1061 2401 -993 2435
rect -903 2401 -835 2435
rect -745 2401 -677 2435
rect -587 2401 -519 2435
rect -429 2401 -361 2435
rect -271 2401 -203 2435
rect -113 2401 -45 2435
rect 45 2401 113 2435
rect 203 2401 271 2435
rect 361 2401 429 2435
rect 519 2401 587 2435
rect 677 2401 745 2435
rect 835 2401 903 2435
rect 993 2401 1061 2435
rect 1151 2401 1219 2435
rect 1309 2401 1377 2435
rect 1467 2401 1535 2435
rect 1625 2401 1693 2435
rect 1783 2401 1851 2435
rect 1941 2401 2009 2435
rect 2099 2401 2167 2435
rect 2257 2401 2325 2435
rect 2415 2401 2483 2435
rect 2573 2401 2641 2435
rect 2731 2401 2799 2435
rect 2889 2401 2957 2435
rect 3047 2401 3115 2435
rect 3205 2401 3273 2435
rect 3363 2401 3431 2435
rect 3521 2401 3589 2435
rect 3679 2401 3747 2435
rect 3837 2401 3905 2435
rect 3995 2401 4063 2435
rect 4153 2401 4221 2435
rect 4311 2401 4379 2435
rect 4469 2401 4537 2435
rect 4627 2401 4695 2435
rect 4785 2401 4853 2435
rect -4853 1273 -4785 1307
rect -4695 1273 -4627 1307
rect -4537 1273 -4469 1307
rect -4379 1273 -4311 1307
rect -4221 1273 -4153 1307
rect -4063 1273 -3995 1307
rect -3905 1273 -3837 1307
rect -3747 1273 -3679 1307
rect -3589 1273 -3521 1307
rect -3431 1273 -3363 1307
rect -3273 1273 -3205 1307
rect -3115 1273 -3047 1307
rect -2957 1273 -2889 1307
rect -2799 1273 -2731 1307
rect -2641 1273 -2573 1307
rect -2483 1273 -2415 1307
rect -2325 1273 -2257 1307
rect -2167 1273 -2099 1307
rect -2009 1273 -1941 1307
rect -1851 1273 -1783 1307
rect -1693 1273 -1625 1307
rect -1535 1273 -1467 1307
rect -1377 1273 -1309 1307
rect -1219 1273 -1151 1307
rect -1061 1273 -993 1307
rect -903 1273 -835 1307
rect -745 1273 -677 1307
rect -587 1273 -519 1307
rect -429 1273 -361 1307
rect -271 1273 -203 1307
rect -113 1273 -45 1307
rect 45 1273 113 1307
rect 203 1273 271 1307
rect 361 1273 429 1307
rect 519 1273 587 1307
rect 677 1273 745 1307
rect 835 1273 903 1307
rect 993 1273 1061 1307
rect 1151 1273 1219 1307
rect 1309 1273 1377 1307
rect 1467 1273 1535 1307
rect 1625 1273 1693 1307
rect 1783 1273 1851 1307
rect 1941 1273 2009 1307
rect 2099 1273 2167 1307
rect 2257 1273 2325 1307
rect 2415 1273 2483 1307
rect 2573 1273 2641 1307
rect 2731 1273 2799 1307
rect 2889 1273 2957 1307
rect 3047 1273 3115 1307
rect 3205 1273 3273 1307
rect 3363 1273 3431 1307
rect 3521 1273 3589 1307
rect 3679 1273 3747 1307
rect 3837 1273 3905 1307
rect 3995 1273 4063 1307
rect 4153 1273 4221 1307
rect 4311 1273 4379 1307
rect 4469 1273 4537 1307
rect 4627 1273 4695 1307
rect 4785 1273 4853 1307
rect -4853 1165 -4785 1199
rect -4695 1165 -4627 1199
rect -4537 1165 -4469 1199
rect -4379 1165 -4311 1199
rect -4221 1165 -4153 1199
rect -4063 1165 -3995 1199
rect -3905 1165 -3837 1199
rect -3747 1165 -3679 1199
rect -3589 1165 -3521 1199
rect -3431 1165 -3363 1199
rect -3273 1165 -3205 1199
rect -3115 1165 -3047 1199
rect -2957 1165 -2889 1199
rect -2799 1165 -2731 1199
rect -2641 1165 -2573 1199
rect -2483 1165 -2415 1199
rect -2325 1165 -2257 1199
rect -2167 1165 -2099 1199
rect -2009 1165 -1941 1199
rect -1851 1165 -1783 1199
rect -1693 1165 -1625 1199
rect -1535 1165 -1467 1199
rect -1377 1165 -1309 1199
rect -1219 1165 -1151 1199
rect -1061 1165 -993 1199
rect -903 1165 -835 1199
rect -745 1165 -677 1199
rect -587 1165 -519 1199
rect -429 1165 -361 1199
rect -271 1165 -203 1199
rect -113 1165 -45 1199
rect 45 1165 113 1199
rect 203 1165 271 1199
rect 361 1165 429 1199
rect 519 1165 587 1199
rect 677 1165 745 1199
rect 835 1165 903 1199
rect 993 1165 1061 1199
rect 1151 1165 1219 1199
rect 1309 1165 1377 1199
rect 1467 1165 1535 1199
rect 1625 1165 1693 1199
rect 1783 1165 1851 1199
rect 1941 1165 2009 1199
rect 2099 1165 2167 1199
rect 2257 1165 2325 1199
rect 2415 1165 2483 1199
rect 2573 1165 2641 1199
rect 2731 1165 2799 1199
rect 2889 1165 2957 1199
rect 3047 1165 3115 1199
rect 3205 1165 3273 1199
rect 3363 1165 3431 1199
rect 3521 1165 3589 1199
rect 3679 1165 3747 1199
rect 3837 1165 3905 1199
rect 3995 1165 4063 1199
rect 4153 1165 4221 1199
rect 4311 1165 4379 1199
rect 4469 1165 4537 1199
rect 4627 1165 4695 1199
rect 4785 1165 4853 1199
rect -4853 37 -4785 71
rect -4695 37 -4627 71
rect -4537 37 -4469 71
rect -4379 37 -4311 71
rect -4221 37 -4153 71
rect -4063 37 -3995 71
rect -3905 37 -3837 71
rect -3747 37 -3679 71
rect -3589 37 -3521 71
rect -3431 37 -3363 71
rect -3273 37 -3205 71
rect -3115 37 -3047 71
rect -2957 37 -2889 71
rect -2799 37 -2731 71
rect -2641 37 -2573 71
rect -2483 37 -2415 71
rect -2325 37 -2257 71
rect -2167 37 -2099 71
rect -2009 37 -1941 71
rect -1851 37 -1783 71
rect -1693 37 -1625 71
rect -1535 37 -1467 71
rect -1377 37 -1309 71
rect -1219 37 -1151 71
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect 1151 37 1219 71
rect 1309 37 1377 71
rect 1467 37 1535 71
rect 1625 37 1693 71
rect 1783 37 1851 71
rect 1941 37 2009 71
rect 2099 37 2167 71
rect 2257 37 2325 71
rect 2415 37 2483 71
rect 2573 37 2641 71
rect 2731 37 2799 71
rect 2889 37 2957 71
rect 3047 37 3115 71
rect 3205 37 3273 71
rect 3363 37 3431 71
rect 3521 37 3589 71
rect 3679 37 3747 71
rect 3837 37 3905 71
rect 3995 37 4063 71
rect 4153 37 4221 71
rect 4311 37 4379 71
rect 4469 37 4537 71
rect 4627 37 4695 71
rect 4785 37 4853 71
rect -4853 -71 -4785 -37
rect -4695 -71 -4627 -37
rect -4537 -71 -4469 -37
rect -4379 -71 -4311 -37
rect -4221 -71 -4153 -37
rect -4063 -71 -3995 -37
rect -3905 -71 -3837 -37
rect -3747 -71 -3679 -37
rect -3589 -71 -3521 -37
rect -3431 -71 -3363 -37
rect -3273 -71 -3205 -37
rect -3115 -71 -3047 -37
rect -2957 -71 -2889 -37
rect -2799 -71 -2731 -37
rect -2641 -71 -2573 -37
rect -2483 -71 -2415 -37
rect -2325 -71 -2257 -37
rect -2167 -71 -2099 -37
rect -2009 -71 -1941 -37
rect -1851 -71 -1783 -37
rect -1693 -71 -1625 -37
rect -1535 -71 -1467 -37
rect -1377 -71 -1309 -37
rect -1219 -71 -1151 -37
rect -1061 -71 -993 -37
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect 993 -71 1061 -37
rect 1151 -71 1219 -37
rect 1309 -71 1377 -37
rect 1467 -71 1535 -37
rect 1625 -71 1693 -37
rect 1783 -71 1851 -37
rect 1941 -71 2009 -37
rect 2099 -71 2167 -37
rect 2257 -71 2325 -37
rect 2415 -71 2483 -37
rect 2573 -71 2641 -37
rect 2731 -71 2799 -37
rect 2889 -71 2957 -37
rect 3047 -71 3115 -37
rect 3205 -71 3273 -37
rect 3363 -71 3431 -37
rect 3521 -71 3589 -37
rect 3679 -71 3747 -37
rect 3837 -71 3905 -37
rect 3995 -71 4063 -37
rect 4153 -71 4221 -37
rect 4311 -71 4379 -37
rect 4469 -71 4537 -37
rect 4627 -71 4695 -37
rect 4785 -71 4853 -37
rect -4853 -1199 -4785 -1165
rect -4695 -1199 -4627 -1165
rect -4537 -1199 -4469 -1165
rect -4379 -1199 -4311 -1165
rect -4221 -1199 -4153 -1165
rect -4063 -1199 -3995 -1165
rect -3905 -1199 -3837 -1165
rect -3747 -1199 -3679 -1165
rect -3589 -1199 -3521 -1165
rect -3431 -1199 -3363 -1165
rect -3273 -1199 -3205 -1165
rect -3115 -1199 -3047 -1165
rect -2957 -1199 -2889 -1165
rect -2799 -1199 -2731 -1165
rect -2641 -1199 -2573 -1165
rect -2483 -1199 -2415 -1165
rect -2325 -1199 -2257 -1165
rect -2167 -1199 -2099 -1165
rect -2009 -1199 -1941 -1165
rect -1851 -1199 -1783 -1165
rect -1693 -1199 -1625 -1165
rect -1535 -1199 -1467 -1165
rect -1377 -1199 -1309 -1165
rect -1219 -1199 -1151 -1165
rect -1061 -1199 -993 -1165
rect -903 -1199 -835 -1165
rect -745 -1199 -677 -1165
rect -587 -1199 -519 -1165
rect -429 -1199 -361 -1165
rect -271 -1199 -203 -1165
rect -113 -1199 -45 -1165
rect 45 -1199 113 -1165
rect 203 -1199 271 -1165
rect 361 -1199 429 -1165
rect 519 -1199 587 -1165
rect 677 -1199 745 -1165
rect 835 -1199 903 -1165
rect 993 -1199 1061 -1165
rect 1151 -1199 1219 -1165
rect 1309 -1199 1377 -1165
rect 1467 -1199 1535 -1165
rect 1625 -1199 1693 -1165
rect 1783 -1199 1851 -1165
rect 1941 -1199 2009 -1165
rect 2099 -1199 2167 -1165
rect 2257 -1199 2325 -1165
rect 2415 -1199 2483 -1165
rect 2573 -1199 2641 -1165
rect 2731 -1199 2799 -1165
rect 2889 -1199 2957 -1165
rect 3047 -1199 3115 -1165
rect 3205 -1199 3273 -1165
rect 3363 -1199 3431 -1165
rect 3521 -1199 3589 -1165
rect 3679 -1199 3747 -1165
rect 3837 -1199 3905 -1165
rect 3995 -1199 4063 -1165
rect 4153 -1199 4221 -1165
rect 4311 -1199 4379 -1165
rect 4469 -1199 4537 -1165
rect 4627 -1199 4695 -1165
rect 4785 -1199 4853 -1165
rect -4853 -1307 -4785 -1273
rect -4695 -1307 -4627 -1273
rect -4537 -1307 -4469 -1273
rect -4379 -1307 -4311 -1273
rect -4221 -1307 -4153 -1273
rect -4063 -1307 -3995 -1273
rect -3905 -1307 -3837 -1273
rect -3747 -1307 -3679 -1273
rect -3589 -1307 -3521 -1273
rect -3431 -1307 -3363 -1273
rect -3273 -1307 -3205 -1273
rect -3115 -1307 -3047 -1273
rect -2957 -1307 -2889 -1273
rect -2799 -1307 -2731 -1273
rect -2641 -1307 -2573 -1273
rect -2483 -1307 -2415 -1273
rect -2325 -1307 -2257 -1273
rect -2167 -1307 -2099 -1273
rect -2009 -1307 -1941 -1273
rect -1851 -1307 -1783 -1273
rect -1693 -1307 -1625 -1273
rect -1535 -1307 -1467 -1273
rect -1377 -1307 -1309 -1273
rect -1219 -1307 -1151 -1273
rect -1061 -1307 -993 -1273
rect -903 -1307 -835 -1273
rect -745 -1307 -677 -1273
rect -587 -1307 -519 -1273
rect -429 -1307 -361 -1273
rect -271 -1307 -203 -1273
rect -113 -1307 -45 -1273
rect 45 -1307 113 -1273
rect 203 -1307 271 -1273
rect 361 -1307 429 -1273
rect 519 -1307 587 -1273
rect 677 -1307 745 -1273
rect 835 -1307 903 -1273
rect 993 -1307 1061 -1273
rect 1151 -1307 1219 -1273
rect 1309 -1307 1377 -1273
rect 1467 -1307 1535 -1273
rect 1625 -1307 1693 -1273
rect 1783 -1307 1851 -1273
rect 1941 -1307 2009 -1273
rect 2099 -1307 2167 -1273
rect 2257 -1307 2325 -1273
rect 2415 -1307 2483 -1273
rect 2573 -1307 2641 -1273
rect 2731 -1307 2799 -1273
rect 2889 -1307 2957 -1273
rect 3047 -1307 3115 -1273
rect 3205 -1307 3273 -1273
rect 3363 -1307 3431 -1273
rect 3521 -1307 3589 -1273
rect 3679 -1307 3747 -1273
rect 3837 -1307 3905 -1273
rect 3995 -1307 4063 -1273
rect 4153 -1307 4221 -1273
rect 4311 -1307 4379 -1273
rect 4469 -1307 4537 -1273
rect 4627 -1307 4695 -1273
rect 4785 -1307 4853 -1273
rect -4853 -2435 -4785 -2401
rect -4695 -2435 -4627 -2401
rect -4537 -2435 -4469 -2401
rect -4379 -2435 -4311 -2401
rect -4221 -2435 -4153 -2401
rect -4063 -2435 -3995 -2401
rect -3905 -2435 -3837 -2401
rect -3747 -2435 -3679 -2401
rect -3589 -2435 -3521 -2401
rect -3431 -2435 -3363 -2401
rect -3273 -2435 -3205 -2401
rect -3115 -2435 -3047 -2401
rect -2957 -2435 -2889 -2401
rect -2799 -2435 -2731 -2401
rect -2641 -2435 -2573 -2401
rect -2483 -2435 -2415 -2401
rect -2325 -2435 -2257 -2401
rect -2167 -2435 -2099 -2401
rect -2009 -2435 -1941 -2401
rect -1851 -2435 -1783 -2401
rect -1693 -2435 -1625 -2401
rect -1535 -2435 -1467 -2401
rect -1377 -2435 -1309 -2401
rect -1219 -2435 -1151 -2401
rect -1061 -2435 -993 -2401
rect -903 -2435 -835 -2401
rect -745 -2435 -677 -2401
rect -587 -2435 -519 -2401
rect -429 -2435 -361 -2401
rect -271 -2435 -203 -2401
rect -113 -2435 -45 -2401
rect 45 -2435 113 -2401
rect 203 -2435 271 -2401
rect 361 -2435 429 -2401
rect 519 -2435 587 -2401
rect 677 -2435 745 -2401
rect 835 -2435 903 -2401
rect 993 -2435 1061 -2401
rect 1151 -2435 1219 -2401
rect 1309 -2435 1377 -2401
rect 1467 -2435 1535 -2401
rect 1625 -2435 1693 -2401
rect 1783 -2435 1851 -2401
rect 1941 -2435 2009 -2401
rect 2099 -2435 2167 -2401
rect 2257 -2435 2325 -2401
rect 2415 -2435 2483 -2401
rect 2573 -2435 2641 -2401
rect 2731 -2435 2799 -2401
rect 2889 -2435 2957 -2401
rect 3047 -2435 3115 -2401
rect 3205 -2435 3273 -2401
rect 3363 -2435 3431 -2401
rect 3521 -2435 3589 -2401
rect 3679 -2435 3747 -2401
rect 3837 -2435 3905 -2401
rect 3995 -2435 4063 -2401
rect 4153 -2435 4221 -2401
rect 4311 -2435 4379 -2401
rect 4469 -2435 4537 -2401
rect 4627 -2435 4695 -2401
rect 4785 -2435 4853 -2401
<< locali >>
rect -5049 2539 -4953 2573
rect 4953 2539 5049 2573
rect -5049 2477 -5015 2539
rect 5015 2477 5049 2539
rect -4869 2401 -4853 2435
rect -4785 2401 -4769 2435
rect -4711 2401 -4695 2435
rect -4627 2401 -4611 2435
rect -4553 2401 -4537 2435
rect -4469 2401 -4453 2435
rect -4395 2401 -4379 2435
rect -4311 2401 -4295 2435
rect -4237 2401 -4221 2435
rect -4153 2401 -4137 2435
rect -4079 2401 -4063 2435
rect -3995 2401 -3979 2435
rect -3921 2401 -3905 2435
rect -3837 2401 -3821 2435
rect -3763 2401 -3747 2435
rect -3679 2401 -3663 2435
rect -3605 2401 -3589 2435
rect -3521 2401 -3505 2435
rect -3447 2401 -3431 2435
rect -3363 2401 -3347 2435
rect -3289 2401 -3273 2435
rect -3205 2401 -3189 2435
rect -3131 2401 -3115 2435
rect -3047 2401 -3031 2435
rect -2973 2401 -2957 2435
rect -2889 2401 -2873 2435
rect -2815 2401 -2799 2435
rect -2731 2401 -2715 2435
rect -2657 2401 -2641 2435
rect -2573 2401 -2557 2435
rect -2499 2401 -2483 2435
rect -2415 2401 -2399 2435
rect -2341 2401 -2325 2435
rect -2257 2401 -2241 2435
rect -2183 2401 -2167 2435
rect -2099 2401 -2083 2435
rect -2025 2401 -2009 2435
rect -1941 2401 -1925 2435
rect -1867 2401 -1851 2435
rect -1783 2401 -1767 2435
rect -1709 2401 -1693 2435
rect -1625 2401 -1609 2435
rect -1551 2401 -1535 2435
rect -1467 2401 -1451 2435
rect -1393 2401 -1377 2435
rect -1309 2401 -1293 2435
rect -1235 2401 -1219 2435
rect -1151 2401 -1135 2435
rect -1077 2401 -1061 2435
rect -993 2401 -977 2435
rect -919 2401 -903 2435
rect -835 2401 -819 2435
rect -761 2401 -745 2435
rect -677 2401 -661 2435
rect -603 2401 -587 2435
rect -519 2401 -503 2435
rect -445 2401 -429 2435
rect -361 2401 -345 2435
rect -287 2401 -271 2435
rect -203 2401 -187 2435
rect -129 2401 -113 2435
rect -45 2401 -29 2435
rect 29 2401 45 2435
rect 113 2401 129 2435
rect 187 2401 203 2435
rect 271 2401 287 2435
rect 345 2401 361 2435
rect 429 2401 445 2435
rect 503 2401 519 2435
rect 587 2401 603 2435
rect 661 2401 677 2435
rect 745 2401 761 2435
rect 819 2401 835 2435
rect 903 2401 919 2435
rect 977 2401 993 2435
rect 1061 2401 1077 2435
rect 1135 2401 1151 2435
rect 1219 2401 1235 2435
rect 1293 2401 1309 2435
rect 1377 2401 1393 2435
rect 1451 2401 1467 2435
rect 1535 2401 1551 2435
rect 1609 2401 1625 2435
rect 1693 2401 1709 2435
rect 1767 2401 1783 2435
rect 1851 2401 1867 2435
rect 1925 2401 1941 2435
rect 2009 2401 2025 2435
rect 2083 2401 2099 2435
rect 2167 2401 2183 2435
rect 2241 2401 2257 2435
rect 2325 2401 2341 2435
rect 2399 2401 2415 2435
rect 2483 2401 2499 2435
rect 2557 2401 2573 2435
rect 2641 2401 2657 2435
rect 2715 2401 2731 2435
rect 2799 2401 2815 2435
rect 2873 2401 2889 2435
rect 2957 2401 2973 2435
rect 3031 2401 3047 2435
rect 3115 2401 3131 2435
rect 3189 2401 3205 2435
rect 3273 2401 3289 2435
rect 3347 2401 3363 2435
rect 3431 2401 3447 2435
rect 3505 2401 3521 2435
rect 3589 2401 3605 2435
rect 3663 2401 3679 2435
rect 3747 2401 3763 2435
rect 3821 2401 3837 2435
rect 3905 2401 3921 2435
rect 3979 2401 3995 2435
rect 4063 2401 4079 2435
rect 4137 2401 4153 2435
rect 4221 2401 4237 2435
rect 4295 2401 4311 2435
rect 4379 2401 4395 2435
rect 4453 2401 4469 2435
rect 4537 2401 4553 2435
rect 4611 2401 4627 2435
rect 4695 2401 4711 2435
rect 4769 2401 4785 2435
rect 4853 2401 4869 2435
rect -4915 2342 -4881 2358
rect -4915 1350 -4881 1366
rect -4757 2342 -4723 2358
rect -4757 1350 -4723 1366
rect -4599 2342 -4565 2358
rect -4599 1350 -4565 1366
rect -4441 2342 -4407 2358
rect -4441 1350 -4407 1366
rect -4283 2342 -4249 2358
rect -4283 1350 -4249 1366
rect -4125 2342 -4091 2358
rect -4125 1350 -4091 1366
rect -3967 2342 -3933 2358
rect -3967 1350 -3933 1366
rect -3809 2342 -3775 2358
rect -3809 1350 -3775 1366
rect -3651 2342 -3617 2358
rect -3651 1350 -3617 1366
rect -3493 2342 -3459 2358
rect -3493 1350 -3459 1366
rect -3335 2342 -3301 2358
rect -3335 1350 -3301 1366
rect -3177 2342 -3143 2358
rect -3177 1350 -3143 1366
rect -3019 2342 -2985 2358
rect -3019 1350 -2985 1366
rect -2861 2342 -2827 2358
rect -2861 1350 -2827 1366
rect -2703 2342 -2669 2358
rect -2703 1350 -2669 1366
rect -2545 2342 -2511 2358
rect -2545 1350 -2511 1366
rect -2387 2342 -2353 2358
rect -2387 1350 -2353 1366
rect -2229 2342 -2195 2358
rect -2229 1350 -2195 1366
rect -2071 2342 -2037 2358
rect -2071 1350 -2037 1366
rect -1913 2342 -1879 2358
rect -1913 1350 -1879 1366
rect -1755 2342 -1721 2358
rect -1755 1350 -1721 1366
rect -1597 2342 -1563 2358
rect -1597 1350 -1563 1366
rect -1439 2342 -1405 2358
rect -1439 1350 -1405 1366
rect -1281 2342 -1247 2358
rect -1281 1350 -1247 1366
rect -1123 2342 -1089 2358
rect -1123 1350 -1089 1366
rect -965 2342 -931 2358
rect -965 1350 -931 1366
rect -807 2342 -773 2358
rect -807 1350 -773 1366
rect -649 2342 -615 2358
rect -649 1350 -615 1366
rect -491 2342 -457 2358
rect -491 1350 -457 1366
rect -333 2342 -299 2358
rect -333 1350 -299 1366
rect -175 2342 -141 2358
rect -175 1350 -141 1366
rect -17 2342 17 2358
rect -17 1350 17 1366
rect 141 2342 175 2358
rect 141 1350 175 1366
rect 299 2342 333 2358
rect 299 1350 333 1366
rect 457 2342 491 2358
rect 457 1350 491 1366
rect 615 2342 649 2358
rect 615 1350 649 1366
rect 773 2342 807 2358
rect 773 1350 807 1366
rect 931 2342 965 2358
rect 931 1350 965 1366
rect 1089 2342 1123 2358
rect 1089 1350 1123 1366
rect 1247 2342 1281 2358
rect 1247 1350 1281 1366
rect 1405 2342 1439 2358
rect 1405 1350 1439 1366
rect 1563 2342 1597 2358
rect 1563 1350 1597 1366
rect 1721 2342 1755 2358
rect 1721 1350 1755 1366
rect 1879 2342 1913 2358
rect 1879 1350 1913 1366
rect 2037 2342 2071 2358
rect 2037 1350 2071 1366
rect 2195 2342 2229 2358
rect 2195 1350 2229 1366
rect 2353 2342 2387 2358
rect 2353 1350 2387 1366
rect 2511 2342 2545 2358
rect 2511 1350 2545 1366
rect 2669 2342 2703 2358
rect 2669 1350 2703 1366
rect 2827 2342 2861 2358
rect 2827 1350 2861 1366
rect 2985 2342 3019 2358
rect 2985 1350 3019 1366
rect 3143 2342 3177 2358
rect 3143 1350 3177 1366
rect 3301 2342 3335 2358
rect 3301 1350 3335 1366
rect 3459 2342 3493 2358
rect 3459 1350 3493 1366
rect 3617 2342 3651 2358
rect 3617 1350 3651 1366
rect 3775 2342 3809 2358
rect 3775 1350 3809 1366
rect 3933 2342 3967 2358
rect 3933 1350 3967 1366
rect 4091 2342 4125 2358
rect 4091 1350 4125 1366
rect 4249 2342 4283 2358
rect 4249 1350 4283 1366
rect 4407 2342 4441 2358
rect 4407 1350 4441 1366
rect 4565 2342 4599 2358
rect 4565 1350 4599 1366
rect 4723 2342 4757 2358
rect 4723 1350 4757 1366
rect 4881 2342 4915 2358
rect 4881 1350 4915 1366
rect -4869 1273 -4853 1307
rect -4785 1273 -4769 1307
rect -4711 1273 -4695 1307
rect -4627 1273 -4611 1307
rect -4553 1273 -4537 1307
rect -4469 1273 -4453 1307
rect -4395 1273 -4379 1307
rect -4311 1273 -4295 1307
rect -4237 1273 -4221 1307
rect -4153 1273 -4137 1307
rect -4079 1273 -4063 1307
rect -3995 1273 -3979 1307
rect -3921 1273 -3905 1307
rect -3837 1273 -3821 1307
rect -3763 1273 -3747 1307
rect -3679 1273 -3663 1307
rect -3605 1273 -3589 1307
rect -3521 1273 -3505 1307
rect -3447 1273 -3431 1307
rect -3363 1273 -3347 1307
rect -3289 1273 -3273 1307
rect -3205 1273 -3189 1307
rect -3131 1273 -3115 1307
rect -3047 1273 -3031 1307
rect -2973 1273 -2957 1307
rect -2889 1273 -2873 1307
rect -2815 1273 -2799 1307
rect -2731 1273 -2715 1307
rect -2657 1273 -2641 1307
rect -2573 1273 -2557 1307
rect -2499 1273 -2483 1307
rect -2415 1273 -2399 1307
rect -2341 1273 -2325 1307
rect -2257 1273 -2241 1307
rect -2183 1273 -2167 1307
rect -2099 1273 -2083 1307
rect -2025 1273 -2009 1307
rect -1941 1273 -1925 1307
rect -1867 1273 -1851 1307
rect -1783 1273 -1767 1307
rect -1709 1273 -1693 1307
rect -1625 1273 -1609 1307
rect -1551 1273 -1535 1307
rect -1467 1273 -1451 1307
rect -1393 1273 -1377 1307
rect -1309 1273 -1293 1307
rect -1235 1273 -1219 1307
rect -1151 1273 -1135 1307
rect -1077 1273 -1061 1307
rect -993 1273 -977 1307
rect -919 1273 -903 1307
rect -835 1273 -819 1307
rect -761 1273 -745 1307
rect -677 1273 -661 1307
rect -603 1273 -587 1307
rect -519 1273 -503 1307
rect -445 1273 -429 1307
rect -361 1273 -345 1307
rect -287 1273 -271 1307
rect -203 1273 -187 1307
rect -129 1273 -113 1307
rect -45 1273 -29 1307
rect 29 1273 45 1307
rect 113 1273 129 1307
rect 187 1273 203 1307
rect 271 1273 287 1307
rect 345 1273 361 1307
rect 429 1273 445 1307
rect 503 1273 519 1307
rect 587 1273 603 1307
rect 661 1273 677 1307
rect 745 1273 761 1307
rect 819 1273 835 1307
rect 903 1273 919 1307
rect 977 1273 993 1307
rect 1061 1273 1077 1307
rect 1135 1273 1151 1307
rect 1219 1273 1235 1307
rect 1293 1273 1309 1307
rect 1377 1273 1393 1307
rect 1451 1273 1467 1307
rect 1535 1273 1551 1307
rect 1609 1273 1625 1307
rect 1693 1273 1709 1307
rect 1767 1273 1783 1307
rect 1851 1273 1867 1307
rect 1925 1273 1941 1307
rect 2009 1273 2025 1307
rect 2083 1273 2099 1307
rect 2167 1273 2183 1307
rect 2241 1273 2257 1307
rect 2325 1273 2341 1307
rect 2399 1273 2415 1307
rect 2483 1273 2499 1307
rect 2557 1273 2573 1307
rect 2641 1273 2657 1307
rect 2715 1273 2731 1307
rect 2799 1273 2815 1307
rect 2873 1273 2889 1307
rect 2957 1273 2973 1307
rect 3031 1273 3047 1307
rect 3115 1273 3131 1307
rect 3189 1273 3205 1307
rect 3273 1273 3289 1307
rect 3347 1273 3363 1307
rect 3431 1273 3447 1307
rect 3505 1273 3521 1307
rect 3589 1273 3605 1307
rect 3663 1273 3679 1307
rect 3747 1273 3763 1307
rect 3821 1273 3837 1307
rect 3905 1273 3921 1307
rect 3979 1273 3995 1307
rect 4063 1273 4079 1307
rect 4137 1273 4153 1307
rect 4221 1273 4237 1307
rect 4295 1273 4311 1307
rect 4379 1273 4395 1307
rect 4453 1273 4469 1307
rect 4537 1273 4553 1307
rect 4611 1273 4627 1307
rect 4695 1273 4711 1307
rect 4769 1273 4785 1307
rect 4853 1273 4869 1307
rect -4869 1165 -4853 1199
rect -4785 1165 -4769 1199
rect -4711 1165 -4695 1199
rect -4627 1165 -4611 1199
rect -4553 1165 -4537 1199
rect -4469 1165 -4453 1199
rect -4395 1165 -4379 1199
rect -4311 1165 -4295 1199
rect -4237 1165 -4221 1199
rect -4153 1165 -4137 1199
rect -4079 1165 -4063 1199
rect -3995 1165 -3979 1199
rect -3921 1165 -3905 1199
rect -3837 1165 -3821 1199
rect -3763 1165 -3747 1199
rect -3679 1165 -3663 1199
rect -3605 1165 -3589 1199
rect -3521 1165 -3505 1199
rect -3447 1165 -3431 1199
rect -3363 1165 -3347 1199
rect -3289 1165 -3273 1199
rect -3205 1165 -3189 1199
rect -3131 1165 -3115 1199
rect -3047 1165 -3031 1199
rect -2973 1165 -2957 1199
rect -2889 1165 -2873 1199
rect -2815 1165 -2799 1199
rect -2731 1165 -2715 1199
rect -2657 1165 -2641 1199
rect -2573 1165 -2557 1199
rect -2499 1165 -2483 1199
rect -2415 1165 -2399 1199
rect -2341 1165 -2325 1199
rect -2257 1165 -2241 1199
rect -2183 1165 -2167 1199
rect -2099 1165 -2083 1199
rect -2025 1165 -2009 1199
rect -1941 1165 -1925 1199
rect -1867 1165 -1851 1199
rect -1783 1165 -1767 1199
rect -1709 1165 -1693 1199
rect -1625 1165 -1609 1199
rect -1551 1165 -1535 1199
rect -1467 1165 -1451 1199
rect -1393 1165 -1377 1199
rect -1309 1165 -1293 1199
rect -1235 1165 -1219 1199
rect -1151 1165 -1135 1199
rect -1077 1165 -1061 1199
rect -993 1165 -977 1199
rect -919 1165 -903 1199
rect -835 1165 -819 1199
rect -761 1165 -745 1199
rect -677 1165 -661 1199
rect -603 1165 -587 1199
rect -519 1165 -503 1199
rect -445 1165 -429 1199
rect -361 1165 -345 1199
rect -287 1165 -271 1199
rect -203 1165 -187 1199
rect -129 1165 -113 1199
rect -45 1165 -29 1199
rect 29 1165 45 1199
rect 113 1165 129 1199
rect 187 1165 203 1199
rect 271 1165 287 1199
rect 345 1165 361 1199
rect 429 1165 445 1199
rect 503 1165 519 1199
rect 587 1165 603 1199
rect 661 1165 677 1199
rect 745 1165 761 1199
rect 819 1165 835 1199
rect 903 1165 919 1199
rect 977 1165 993 1199
rect 1061 1165 1077 1199
rect 1135 1165 1151 1199
rect 1219 1165 1235 1199
rect 1293 1165 1309 1199
rect 1377 1165 1393 1199
rect 1451 1165 1467 1199
rect 1535 1165 1551 1199
rect 1609 1165 1625 1199
rect 1693 1165 1709 1199
rect 1767 1165 1783 1199
rect 1851 1165 1867 1199
rect 1925 1165 1941 1199
rect 2009 1165 2025 1199
rect 2083 1165 2099 1199
rect 2167 1165 2183 1199
rect 2241 1165 2257 1199
rect 2325 1165 2341 1199
rect 2399 1165 2415 1199
rect 2483 1165 2499 1199
rect 2557 1165 2573 1199
rect 2641 1165 2657 1199
rect 2715 1165 2731 1199
rect 2799 1165 2815 1199
rect 2873 1165 2889 1199
rect 2957 1165 2973 1199
rect 3031 1165 3047 1199
rect 3115 1165 3131 1199
rect 3189 1165 3205 1199
rect 3273 1165 3289 1199
rect 3347 1165 3363 1199
rect 3431 1165 3447 1199
rect 3505 1165 3521 1199
rect 3589 1165 3605 1199
rect 3663 1165 3679 1199
rect 3747 1165 3763 1199
rect 3821 1165 3837 1199
rect 3905 1165 3921 1199
rect 3979 1165 3995 1199
rect 4063 1165 4079 1199
rect 4137 1165 4153 1199
rect 4221 1165 4237 1199
rect 4295 1165 4311 1199
rect 4379 1165 4395 1199
rect 4453 1165 4469 1199
rect 4537 1165 4553 1199
rect 4611 1165 4627 1199
rect 4695 1165 4711 1199
rect 4769 1165 4785 1199
rect 4853 1165 4869 1199
rect -4915 1106 -4881 1122
rect -4915 114 -4881 130
rect -4757 1106 -4723 1122
rect -4757 114 -4723 130
rect -4599 1106 -4565 1122
rect -4599 114 -4565 130
rect -4441 1106 -4407 1122
rect -4441 114 -4407 130
rect -4283 1106 -4249 1122
rect -4283 114 -4249 130
rect -4125 1106 -4091 1122
rect -4125 114 -4091 130
rect -3967 1106 -3933 1122
rect -3967 114 -3933 130
rect -3809 1106 -3775 1122
rect -3809 114 -3775 130
rect -3651 1106 -3617 1122
rect -3651 114 -3617 130
rect -3493 1106 -3459 1122
rect -3493 114 -3459 130
rect -3335 1106 -3301 1122
rect -3335 114 -3301 130
rect -3177 1106 -3143 1122
rect -3177 114 -3143 130
rect -3019 1106 -2985 1122
rect -3019 114 -2985 130
rect -2861 1106 -2827 1122
rect -2861 114 -2827 130
rect -2703 1106 -2669 1122
rect -2703 114 -2669 130
rect -2545 1106 -2511 1122
rect -2545 114 -2511 130
rect -2387 1106 -2353 1122
rect -2387 114 -2353 130
rect -2229 1106 -2195 1122
rect -2229 114 -2195 130
rect -2071 1106 -2037 1122
rect -2071 114 -2037 130
rect -1913 1106 -1879 1122
rect -1913 114 -1879 130
rect -1755 1106 -1721 1122
rect -1755 114 -1721 130
rect -1597 1106 -1563 1122
rect -1597 114 -1563 130
rect -1439 1106 -1405 1122
rect -1439 114 -1405 130
rect -1281 1106 -1247 1122
rect -1281 114 -1247 130
rect -1123 1106 -1089 1122
rect -1123 114 -1089 130
rect -965 1106 -931 1122
rect -965 114 -931 130
rect -807 1106 -773 1122
rect -807 114 -773 130
rect -649 1106 -615 1122
rect -649 114 -615 130
rect -491 1106 -457 1122
rect -491 114 -457 130
rect -333 1106 -299 1122
rect -333 114 -299 130
rect -175 1106 -141 1122
rect -175 114 -141 130
rect -17 1106 17 1122
rect -17 114 17 130
rect 141 1106 175 1122
rect 141 114 175 130
rect 299 1106 333 1122
rect 299 114 333 130
rect 457 1106 491 1122
rect 457 114 491 130
rect 615 1106 649 1122
rect 615 114 649 130
rect 773 1106 807 1122
rect 773 114 807 130
rect 931 1106 965 1122
rect 931 114 965 130
rect 1089 1106 1123 1122
rect 1089 114 1123 130
rect 1247 1106 1281 1122
rect 1247 114 1281 130
rect 1405 1106 1439 1122
rect 1405 114 1439 130
rect 1563 1106 1597 1122
rect 1563 114 1597 130
rect 1721 1106 1755 1122
rect 1721 114 1755 130
rect 1879 1106 1913 1122
rect 1879 114 1913 130
rect 2037 1106 2071 1122
rect 2037 114 2071 130
rect 2195 1106 2229 1122
rect 2195 114 2229 130
rect 2353 1106 2387 1122
rect 2353 114 2387 130
rect 2511 1106 2545 1122
rect 2511 114 2545 130
rect 2669 1106 2703 1122
rect 2669 114 2703 130
rect 2827 1106 2861 1122
rect 2827 114 2861 130
rect 2985 1106 3019 1122
rect 2985 114 3019 130
rect 3143 1106 3177 1122
rect 3143 114 3177 130
rect 3301 1106 3335 1122
rect 3301 114 3335 130
rect 3459 1106 3493 1122
rect 3459 114 3493 130
rect 3617 1106 3651 1122
rect 3617 114 3651 130
rect 3775 1106 3809 1122
rect 3775 114 3809 130
rect 3933 1106 3967 1122
rect 3933 114 3967 130
rect 4091 1106 4125 1122
rect 4091 114 4125 130
rect 4249 1106 4283 1122
rect 4249 114 4283 130
rect 4407 1106 4441 1122
rect 4407 114 4441 130
rect 4565 1106 4599 1122
rect 4565 114 4599 130
rect 4723 1106 4757 1122
rect 4723 114 4757 130
rect 4881 1106 4915 1122
rect 4881 114 4915 130
rect -4869 37 -4853 71
rect -4785 37 -4769 71
rect -4711 37 -4695 71
rect -4627 37 -4611 71
rect -4553 37 -4537 71
rect -4469 37 -4453 71
rect -4395 37 -4379 71
rect -4311 37 -4295 71
rect -4237 37 -4221 71
rect -4153 37 -4137 71
rect -4079 37 -4063 71
rect -3995 37 -3979 71
rect -3921 37 -3905 71
rect -3837 37 -3821 71
rect -3763 37 -3747 71
rect -3679 37 -3663 71
rect -3605 37 -3589 71
rect -3521 37 -3505 71
rect -3447 37 -3431 71
rect -3363 37 -3347 71
rect -3289 37 -3273 71
rect -3205 37 -3189 71
rect -3131 37 -3115 71
rect -3047 37 -3031 71
rect -2973 37 -2957 71
rect -2889 37 -2873 71
rect -2815 37 -2799 71
rect -2731 37 -2715 71
rect -2657 37 -2641 71
rect -2573 37 -2557 71
rect -2499 37 -2483 71
rect -2415 37 -2399 71
rect -2341 37 -2325 71
rect -2257 37 -2241 71
rect -2183 37 -2167 71
rect -2099 37 -2083 71
rect -2025 37 -2009 71
rect -1941 37 -1925 71
rect -1867 37 -1851 71
rect -1783 37 -1767 71
rect -1709 37 -1693 71
rect -1625 37 -1609 71
rect -1551 37 -1535 71
rect -1467 37 -1451 71
rect -1393 37 -1377 71
rect -1309 37 -1293 71
rect -1235 37 -1219 71
rect -1151 37 -1135 71
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -919 37 -903 71
rect -835 37 -819 71
rect -761 37 -745 71
rect -677 37 -661 71
rect -603 37 -587 71
rect -519 37 -503 71
rect -445 37 -429 71
rect -361 37 -345 71
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect 345 37 361 71
rect 429 37 445 71
rect 503 37 519 71
rect 587 37 603 71
rect 661 37 677 71
rect 745 37 761 71
rect 819 37 835 71
rect 903 37 919 71
rect 977 37 993 71
rect 1061 37 1077 71
rect 1135 37 1151 71
rect 1219 37 1235 71
rect 1293 37 1309 71
rect 1377 37 1393 71
rect 1451 37 1467 71
rect 1535 37 1551 71
rect 1609 37 1625 71
rect 1693 37 1709 71
rect 1767 37 1783 71
rect 1851 37 1867 71
rect 1925 37 1941 71
rect 2009 37 2025 71
rect 2083 37 2099 71
rect 2167 37 2183 71
rect 2241 37 2257 71
rect 2325 37 2341 71
rect 2399 37 2415 71
rect 2483 37 2499 71
rect 2557 37 2573 71
rect 2641 37 2657 71
rect 2715 37 2731 71
rect 2799 37 2815 71
rect 2873 37 2889 71
rect 2957 37 2973 71
rect 3031 37 3047 71
rect 3115 37 3131 71
rect 3189 37 3205 71
rect 3273 37 3289 71
rect 3347 37 3363 71
rect 3431 37 3447 71
rect 3505 37 3521 71
rect 3589 37 3605 71
rect 3663 37 3679 71
rect 3747 37 3763 71
rect 3821 37 3837 71
rect 3905 37 3921 71
rect 3979 37 3995 71
rect 4063 37 4079 71
rect 4137 37 4153 71
rect 4221 37 4237 71
rect 4295 37 4311 71
rect 4379 37 4395 71
rect 4453 37 4469 71
rect 4537 37 4553 71
rect 4611 37 4627 71
rect 4695 37 4711 71
rect 4769 37 4785 71
rect 4853 37 4869 71
rect -4869 -71 -4853 -37
rect -4785 -71 -4769 -37
rect -4711 -71 -4695 -37
rect -4627 -71 -4611 -37
rect -4553 -71 -4537 -37
rect -4469 -71 -4453 -37
rect -4395 -71 -4379 -37
rect -4311 -71 -4295 -37
rect -4237 -71 -4221 -37
rect -4153 -71 -4137 -37
rect -4079 -71 -4063 -37
rect -3995 -71 -3979 -37
rect -3921 -71 -3905 -37
rect -3837 -71 -3821 -37
rect -3763 -71 -3747 -37
rect -3679 -71 -3663 -37
rect -3605 -71 -3589 -37
rect -3521 -71 -3505 -37
rect -3447 -71 -3431 -37
rect -3363 -71 -3347 -37
rect -3289 -71 -3273 -37
rect -3205 -71 -3189 -37
rect -3131 -71 -3115 -37
rect -3047 -71 -3031 -37
rect -2973 -71 -2957 -37
rect -2889 -71 -2873 -37
rect -2815 -71 -2799 -37
rect -2731 -71 -2715 -37
rect -2657 -71 -2641 -37
rect -2573 -71 -2557 -37
rect -2499 -71 -2483 -37
rect -2415 -71 -2399 -37
rect -2341 -71 -2325 -37
rect -2257 -71 -2241 -37
rect -2183 -71 -2167 -37
rect -2099 -71 -2083 -37
rect -2025 -71 -2009 -37
rect -1941 -71 -1925 -37
rect -1867 -71 -1851 -37
rect -1783 -71 -1767 -37
rect -1709 -71 -1693 -37
rect -1625 -71 -1609 -37
rect -1551 -71 -1535 -37
rect -1467 -71 -1451 -37
rect -1393 -71 -1377 -37
rect -1309 -71 -1293 -37
rect -1235 -71 -1219 -37
rect -1151 -71 -1135 -37
rect -1077 -71 -1061 -37
rect -993 -71 -977 -37
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 977 -71 993 -37
rect 1061 -71 1077 -37
rect 1135 -71 1151 -37
rect 1219 -71 1235 -37
rect 1293 -71 1309 -37
rect 1377 -71 1393 -37
rect 1451 -71 1467 -37
rect 1535 -71 1551 -37
rect 1609 -71 1625 -37
rect 1693 -71 1709 -37
rect 1767 -71 1783 -37
rect 1851 -71 1867 -37
rect 1925 -71 1941 -37
rect 2009 -71 2025 -37
rect 2083 -71 2099 -37
rect 2167 -71 2183 -37
rect 2241 -71 2257 -37
rect 2325 -71 2341 -37
rect 2399 -71 2415 -37
rect 2483 -71 2499 -37
rect 2557 -71 2573 -37
rect 2641 -71 2657 -37
rect 2715 -71 2731 -37
rect 2799 -71 2815 -37
rect 2873 -71 2889 -37
rect 2957 -71 2973 -37
rect 3031 -71 3047 -37
rect 3115 -71 3131 -37
rect 3189 -71 3205 -37
rect 3273 -71 3289 -37
rect 3347 -71 3363 -37
rect 3431 -71 3447 -37
rect 3505 -71 3521 -37
rect 3589 -71 3605 -37
rect 3663 -71 3679 -37
rect 3747 -71 3763 -37
rect 3821 -71 3837 -37
rect 3905 -71 3921 -37
rect 3979 -71 3995 -37
rect 4063 -71 4079 -37
rect 4137 -71 4153 -37
rect 4221 -71 4237 -37
rect 4295 -71 4311 -37
rect 4379 -71 4395 -37
rect 4453 -71 4469 -37
rect 4537 -71 4553 -37
rect 4611 -71 4627 -37
rect 4695 -71 4711 -37
rect 4769 -71 4785 -37
rect 4853 -71 4869 -37
rect -4915 -130 -4881 -114
rect -4915 -1122 -4881 -1106
rect -4757 -130 -4723 -114
rect -4757 -1122 -4723 -1106
rect -4599 -130 -4565 -114
rect -4599 -1122 -4565 -1106
rect -4441 -130 -4407 -114
rect -4441 -1122 -4407 -1106
rect -4283 -130 -4249 -114
rect -4283 -1122 -4249 -1106
rect -4125 -130 -4091 -114
rect -4125 -1122 -4091 -1106
rect -3967 -130 -3933 -114
rect -3967 -1122 -3933 -1106
rect -3809 -130 -3775 -114
rect -3809 -1122 -3775 -1106
rect -3651 -130 -3617 -114
rect -3651 -1122 -3617 -1106
rect -3493 -130 -3459 -114
rect -3493 -1122 -3459 -1106
rect -3335 -130 -3301 -114
rect -3335 -1122 -3301 -1106
rect -3177 -130 -3143 -114
rect -3177 -1122 -3143 -1106
rect -3019 -130 -2985 -114
rect -3019 -1122 -2985 -1106
rect -2861 -130 -2827 -114
rect -2861 -1122 -2827 -1106
rect -2703 -130 -2669 -114
rect -2703 -1122 -2669 -1106
rect -2545 -130 -2511 -114
rect -2545 -1122 -2511 -1106
rect -2387 -130 -2353 -114
rect -2387 -1122 -2353 -1106
rect -2229 -130 -2195 -114
rect -2229 -1122 -2195 -1106
rect -2071 -130 -2037 -114
rect -2071 -1122 -2037 -1106
rect -1913 -130 -1879 -114
rect -1913 -1122 -1879 -1106
rect -1755 -130 -1721 -114
rect -1755 -1122 -1721 -1106
rect -1597 -130 -1563 -114
rect -1597 -1122 -1563 -1106
rect -1439 -130 -1405 -114
rect -1439 -1122 -1405 -1106
rect -1281 -130 -1247 -114
rect -1281 -1122 -1247 -1106
rect -1123 -130 -1089 -114
rect -1123 -1122 -1089 -1106
rect -965 -130 -931 -114
rect -965 -1122 -931 -1106
rect -807 -130 -773 -114
rect -807 -1122 -773 -1106
rect -649 -130 -615 -114
rect -649 -1122 -615 -1106
rect -491 -130 -457 -114
rect -491 -1122 -457 -1106
rect -333 -130 -299 -114
rect -333 -1122 -299 -1106
rect -175 -130 -141 -114
rect -175 -1122 -141 -1106
rect -17 -130 17 -114
rect -17 -1122 17 -1106
rect 141 -130 175 -114
rect 141 -1122 175 -1106
rect 299 -130 333 -114
rect 299 -1122 333 -1106
rect 457 -130 491 -114
rect 457 -1122 491 -1106
rect 615 -130 649 -114
rect 615 -1122 649 -1106
rect 773 -130 807 -114
rect 773 -1122 807 -1106
rect 931 -130 965 -114
rect 931 -1122 965 -1106
rect 1089 -130 1123 -114
rect 1089 -1122 1123 -1106
rect 1247 -130 1281 -114
rect 1247 -1122 1281 -1106
rect 1405 -130 1439 -114
rect 1405 -1122 1439 -1106
rect 1563 -130 1597 -114
rect 1563 -1122 1597 -1106
rect 1721 -130 1755 -114
rect 1721 -1122 1755 -1106
rect 1879 -130 1913 -114
rect 1879 -1122 1913 -1106
rect 2037 -130 2071 -114
rect 2037 -1122 2071 -1106
rect 2195 -130 2229 -114
rect 2195 -1122 2229 -1106
rect 2353 -130 2387 -114
rect 2353 -1122 2387 -1106
rect 2511 -130 2545 -114
rect 2511 -1122 2545 -1106
rect 2669 -130 2703 -114
rect 2669 -1122 2703 -1106
rect 2827 -130 2861 -114
rect 2827 -1122 2861 -1106
rect 2985 -130 3019 -114
rect 2985 -1122 3019 -1106
rect 3143 -130 3177 -114
rect 3143 -1122 3177 -1106
rect 3301 -130 3335 -114
rect 3301 -1122 3335 -1106
rect 3459 -130 3493 -114
rect 3459 -1122 3493 -1106
rect 3617 -130 3651 -114
rect 3617 -1122 3651 -1106
rect 3775 -130 3809 -114
rect 3775 -1122 3809 -1106
rect 3933 -130 3967 -114
rect 3933 -1122 3967 -1106
rect 4091 -130 4125 -114
rect 4091 -1122 4125 -1106
rect 4249 -130 4283 -114
rect 4249 -1122 4283 -1106
rect 4407 -130 4441 -114
rect 4407 -1122 4441 -1106
rect 4565 -130 4599 -114
rect 4565 -1122 4599 -1106
rect 4723 -130 4757 -114
rect 4723 -1122 4757 -1106
rect 4881 -130 4915 -114
rect 4881 -1122 4915 -1106
rect -4869 -1199 -4853 -1165
rect -4785 -1199 -4769 -1165
rect -4711 -1199 -4695 -1165
rect -4627 -1199 -4611 -1165
rect -4553 -1199 -4537 -1165
rect -4469 -1199 -4453 -1165
rect -4395 -1199 -4379 -1165
rect -4311 -1199 -4295 -1165
rect -4237 -1199 -4221 -1165
rect -4153 -1199 -4137 -1165
rect -4079 -1199 -4063 -1165
rect -3995 -1199 -3979 -1165
rect -3921 -1199 -3905 -1165
rect -3837 -1199 -3821 -1165
rect -3763 -1199 -3747 -1165
rect -3679 -1199 -3663 -1165
rect -3605 -1199 -3589 -1165
rect -3521 -1199 -3505 -1165
rect -3447 -1199 -3431 -1165
rect -3363 -1199 -3347 -1165
rect -3289 -1199 -3273 -1165
rect -3205 -1199 -3189 -1165
rect -3131 -1199 -3115 -1165
rect -3047 -1199 -3031 -1165
rect -2973 -1199 -2957 -1165
rect -2889 -1199 -2873 -1165
rect -2815 -1199 -2799 -1165
rect -2731 -1199 -2715 -1165
rect -2657 -1199 -2641 -1165
rect -2573 -1199 -2557 -1165
rect -2499 -1199 -2483 -1165
rect -2415 -1199 -2399 -1165
rect -2341 -1199 -2325 -1165
rect -2257 -1199 -2241 -1165
rect -2183 -1199 -2167 -1165
rect -2099 -1199 -2083 -1165
rect -2025 -1199 -2009 -1165
rect -1941 -1199 -1925 -1165
rect -1867 -1199 -1851 -1165
rect -1783 -1199 -1767 -1165
rect -1709 -1199 -1693 -1165
rect -1625 -1199 -1609 -1165
rect -1551 -1199 -1535 -1165
rect -1467 -1199 -1451 -1165
rect -1393 -1199 -1377 -1165
rect -1309 -1199 -1293 -1165
rect -1235 -1199 -1219 -1165
rect -1151 -1199 -1135 -1165
rect -1077 -1199 -1061 -1165
rect -993 -1199 -977 -1165
rect -919 -1199 -903 -1165
rect -835 -1199 -819 -1165
rect -761 -1199 -745 -1165
rect -677 -1199 -661 -1165
rect -603 -1199 -587 -1165
rect -519 -1199 -503 -1165
rect -445 -1199 -429 -1165
rect -361 -1199 -345 -1165
rect -287 -1199 -271 -1165
rect -203 -1199 -187 -1165
rect -129 -1199 -113 -1165
rect -45 -1199 -29 -1165
rect 29 -1199 45 -1165
rect 113 -1199 129 -1165
rect 187 -1199 203 -1165
rect 271 -1199 287 -1165
rect 345 -1199 361 -1165
rect 429 -1199 445 -1165
rect 503 -1199 519 -1165
rect 587 -1199 603 -1165
rect 661 -1199 677 -1165
rect 745 -1199 761 -1165
rect 819 -1199 835 -1165
rect 903 -1199 919 -1165
rect 977 -1199 993 -1165
rect 1061 -1199 1077 -1165
rect 1135 -1199 1151 -1165
rect 1219 -1199 1235 -1165
rect 1293 -1199 1309 -1165
rect 1377 -1199 1393 -1165
rect 1451 -1199 1467 -1165
rect 1535 -1199 1551 -1165
rect 1609 -1199 1625 -1165
rect 1693 -1199 1709 -1165
rect 1767 -1199 1783 -1165
rect 1851 -1199 1867 -1165
rect 1925 -1199 1941 -1165
rect 2009 -1199 2025 -1165
rect 2083 -1199 2099 -1165
rect 2167 -1199 2183 -1165
rect 2241 -1199 2257 -1165
rect 2325 -1199 2341 -1165
rect 2399 -1199 2415 -1165
rect 2483 -1199 2499 -1165
rect 2557 -1199 2573 -1165
rect 2641 -1199 2657 -1165
rect 2715 -1199 2731 -1165
rect 2799 -1199 2815 -1165
rect 2873 -1199 2889 -1165
rect 2957 -1199 2973 -1165
rect 3031 -1199 3047 -1165
rect 3115 -1199 3131 -1165
rect 3189 -1199 3205 -1165
rect 3273 -1199 3289 -1165
rect 3347 -1199 3363 -1165
rect 3431 -1199 3447 -1165
rect 3505 -1199 3521 -1165
rect 3589 -1199 3605 -1165
rect 3663 -1199 3679 -1165
rect 3747 -1199 3763 -1165
rect 3821 -1199 3837 -1165
rect 3905 -1199 3921 -1165
rect 3979 -1199 3995 -1165
rect 4063 -1199 4079 -1165
rect 4137 -1199 4153 -1165
rect 4221 -1199 4237 -1165
rect 4295 -1199 4311 -1165
rect 4379 -1199 4395 -1165
rect 4453 -1199 4469 -1165
rect 4537 -1199 4553 -1165
rect 4611 -1199 4627 -1165
rect 4695 -1199 4711 -1165
rect 4769 -1199 4785 -1165
rect 4853 -1199 4869 -1165
rect -4869 -1307 -4853 -1273
rect -4785 -1307 -4769 -1273
rect -4711 -1307 -4695 -1273
rect -4627 -1307 -4611 -1273
rect -4553 -1307 -4537 -1273
rect -4469 -1307 -4453 -1273
rect -4395 -1307 -4379 -1273
rect -4311 -1307 -4295 -1273
rect -4237 -1307 -4221 -1273
rect -4153 -1307 -4137 -1273
rect -4079 -1307 -4063 -1273
rect -3995 -1307 -3979 -1273
rect -3921 -1307 -3905 -1273
rect -3837 -1307 -3821 -1273
rect -3763 -1307 -3747 -1273
rect -3679 -1307 -3663 -1273
rect -3605 -1307 -3589 -1273
rect -3521 -1307 -3505 -1273
rect -3447 -1307 -3431 -1273
rect -3363 -1307 -3347 -1273
rect -3289 -1307 -3273 -1273
rect -3205 -1307 -3189 -1273
rect -3131 -1307 -3115 -1273
rect -3047 -1307 -3031 -1273
rect -2973 -1307 -2957 -1273
rect -2889 -1307 -2873 -1273
rect -2815 -1307 -2799 -1273
rect -2731 -1307 -2715 -1273
rect -2657 -1307 -2641 -1273
rect -2573 -1307 -2557 -1273
rect -2499 -1307 -2483 -1273
rect -2415 -1307 -2399 -1273
rect -2341 -1307 -2325 -1273
rect -2257 -1307 -2241 -1273
rect -2183 -1307 -2167 -1273
rect -2099 -1307 -2083 -1273
rect -2025 -1307 -2009 -1273
rect -1941 -1307 -1925 -1273
rect -1867 -1307 -1851 -1273
rect -1783 -1307 -1767 -1273
rect -1709 -1307 -1693 -1273
rect -1625 -1307 -1609 -1273
rect -1551 -1307 -1535 -1273
rect -1467 -1307 -1451 -1273
rect -1393 -1307 -1377 -1273
rect -1309 -1307 -1293 -1273
rect -1235 -1307 -1219 -1273
rect -1151 -1307 -1135 -1273
rect -1077 -1307 -1061 -1273
rect -993 -1307 -977 -1273
rect -919 -1307 -903 -1273
rect -835 -1307 -819 -1273
rect -761 -1307 -745 -1273
rect -677 -1307 -661 -1273
rect -603 -1307 -587 -1273
rect -519 -1307 -503 -1273
rect -445 -1307 -429 -1273
rect -361 -1307 -345 -1273
rect -287 -1307 -271 -1273
rect -203 -1307 -187 -1273
rect -129 -1307 -113 -1273
rect -45 -1307 -29 -1273
rect 29 -1307 45 -1273
rect 113 -1307 129 -1273
rect 187 -1307 203 -1273
rect 271 -1307 287 -1273
rect 345 -1307 361 -1273
rect 429 -1307 445 -1273
rect 503 -1307 519 -1273
rect 587 -1307 603 -1273
rect 661 -1307 677 -1273
rect 745 -1307 761 -1273
rect 819 -1307 835 -1273
rect 903 -1307 919 -1273
rect 977 -1307 993 -1273
rect 1061 -1307 1077 -1273
rect 1135 -1307 1151 -1273
rect 1219 -1307 1235 -1273
rect 1293 -1307 1309 -1273
rect 1377 -1307 1393 -1273
rect 1451 -1307 1467 -1273
rect 1535 -1307 1551 -1273
rect 1609 -1307 1625 -1273
rect 1693 -1307 1709 -1273
rect 1767 -1307 1783 -1273
rect 1851 -1307 1867 -1273
rect 1925 -1307 1941 -1273
rect 2009 -1307 2025 -1273
rect 2083 -1307 2099 -1273
rect 2167 -1307 2183 -1273
rect 2241 -1307 2257 -1273
rect 2325 -1307 2341 -1273
rect 2399 -1307 2415 -1273
rect 2483 -1307 2499 -1273
rect 2557 -1307 2573 -1273
rect 2641 -1307 2657 -1273
rect 2715 -1307 2731 -1273
rect 2799 -1307 2815 -1273
rect 2873 -1307 2889 -1273
rect 2957 -1307 2973 -1273
rect 3031 -1307 3047 -1273
rect 3115 -1307 3131 -1273
rect 3189 -1307 3205 -1273
rect 3273 -1307 3289 -1273
rect 3347 -1307 3363 -1273
rect 3431 -1307 3447 -1273
rect 3505 -1307 3521 -1273
rect 3589 -1307 3605 -1273
rect 3663 -1307 3679 -1273
rect 3747 -1307 3763 -1273
rect 3821 -1307 3837 -1273
rect 3905 -1307 3921 -1273
rect 3979 -1307 3995 -1273
rect 4063 -1307 4079 -1273
rect 4137 -1307 4153 -1273
rect 4221 -1307 4237 -1273
rect 4295 -1307 4311 -1273
rect 4379 -1307 4395 -1273
rect 4453 -1307 4469 -1273
rect 4537 -1307 4553 -1273
rect 4611 -1307 4627 -1273
rect 4695 -1307 4711 -1273
rect 4769 -1307 4785 -1273
rect 4853 -1307 4869 -1273
rect -4915 -1366 -4881 -1350
rect -4915 -2358 -4881 -2342
rect -4757 -1366 -4723 -1350
rect -4757 -2358 -4723 -2342
rect -4599 -1366 -4565 -1350
rect -4599 -2358 -4565 -2342
rect -4441 -1366 -4407 -1350
rect -4441 -2358 -4407 -2342
rect -4283 -1366 -4249 -1350
rect -4283 -2358 -4249 -2342
rect -4125 -1366 -4091 -1350
rect -4125 -2358 -4091 -2342
rect -3967 -1366 -3933 -1350
rect -3967 -2358 -3933 -2342
rect -3809 -1366 -3775 -1350
rect -3809 -2358 -3775 -2342
rect -3651 -1366 -3617 -1350
rect -3651 -2358 -3617 -2342
rect -3493 -1366 -3459 -1350
rect -3493 -2358 -3459 -2342
rect -3335 -1366 -3301 -1350
rect -3335 -2358 -3301 -2342
rect -3177 -1366 -3143 -1350
rect -3177 -2358 -3143 -2342
rect -3019 -1366 -2985 -1350
rect -3019 -2358 -2985 -2342
rect -2861 -1366 -2827 -1350
rect -2861 -2358 -2827 -2342
rect -2703 -1366 -2669 -1350
rect -2703 -2358 -2669 -2342
rect -2545 -1366 -2511 -1350
rect -2545 -2358 -2511 -2342
rect -2387 -1366 -2353 -1350
rect -2387 -2358 -2353 -2342
rect -2229 -1366 -2195 -1350
rect -2229 -2358 -2195 -2342
rect -2071 -1366 -2037 -1350
rect -2071 -2358 -2037 -2342
rect -1913 -1366 -1879 -1350
rect -1913 -2358 -1879 -2342
rect -1755 -1366 -1721 -1350
rect -1755 -2358 -1721 -2342
rect -1597 -1366 -1563 -1350
rect -1597 -2358 -1563 -2342
rect -1439 -1366 -1405 -1350
rect -1439 -2358 -1405 -2342
rect -1281 -1366 -1247 -1350
rect -1281 -2358 -1247 -2342
rect -1123 -1366 -1089 -1350
rect -1123 -2358 -1089 -2342
rect -965 -1366 -931 -1350
rect -965 -2358 -931 -2342
rect -807 -1366 -773 -1350
rect -807 -2358 -773 -2342
rect -649 -1366 -615 -1350
rect -649 -2358 -615 -2342
rect -491 -1366 -457 -1350
rect -491 -2358 -457 -2342
rect -333 -1366 -299 -1350
rect -333 -2358 -299 -2342
rect -175 -1366 -141 -1350
rect -175 -2358 -141 -2342
rect -17 -1366 17 -1350
rect -17 -2358 17 -2342
rect 141 -1366 175 -1350
rect 141 -2358 175 -2342
rect 299 -1366 333 -1350
rect 299 -2358 333 -2342
rect 457 -1366 491 -1350
rect 457 -2358 491 -2342
rect 615 -1366 649 -1350
rect 615 -2358 649 -2342
rect 773 -1366 807 -1350
rect 773 -2358 807 -2342
rect 931 -1366 965 -1350
rect 931 -2358 965 -2342
rect 1089 -1366 1123 -1350
rect 1089 -2358 1123 -2342
rect 1247 -1366 1281 -1350
rect 1247 -2358 1281 -2342
rect 1405 -1366 1439 -1350
rect 1405 -2358 1439 -2342
rect 1563 -1366 1597 -1350
rect 1563 -2358 1597 -2342
rect 1721 -1366 1755 -1350
rect 1721 -2358 1755 -2342
rect 1879 -1366 1913 -1350
rect 1879 -2358 1913 -2342
rect 2037 -1366 2071 -1350
rect 2037 -2358 2071 -2342
rect 2195 -1366 2229 -1350
rect 2195 -2358 2229 -2342
rect 2353 -1366 2387 -1350
rect 2353 -2358 2387 -2342
rect 2511 -1366 2545 -1350
rect 2511 -2358 2545 -2342
rect 2669 -1366 2703 -1350
rect 2669 -2358 2703 -2342
rect 2827 -1366 2861 -1350
rect 2827 -2358 2861 -2342
rect 2985 -1366 3019 -1350
rect 2985 -2358 3019 -2342
rect 3143 -1366 3177 -1350
rect 3143 -2358 3177 -2342
rect 3301 -1366 3335 -1350
rect 3301 -2358 3335 -2342
rect 3459 -1366 3493 -1350
rect 3459 -2358 3493 -2342
rect 3617 -1366 3651 -1350
rect 3617 -2358 3651 -2342
rect 3775 -1366 3809 -1350
rect 3775 -2358 3809 -2342
rect 3933 -1366 3967 -1350
rect 3933 -2358 3967 -2342
rect 4091 -1366 4125 -1350
rect 4091 -2358 4125 -2342
rect 4249 -1366 4283 -1350
rect 4249 -2358 4283 -2342
rect 4407 -1366 4441 -1350
rect 4407 -2358 4441 -2342
rect 4565 -1366 4599 -1350
rect 4565 -2358 4599 -2342
rect 4723 -1366 4757 -1350
rect 4723 -2358 4757 -2342
rect 4881 -1366 4915 -1350
rect 4881 -2358 4915 -2342
rect -4869 -2435 -4853 -2401
rect -4785 -2435 -4769 -2401
rect -4711 -2435 -4695 -2401
rect -4627 -2435 -4611 -2401
rect -4553 -2435 -4537 -2401
rect -4469 -2435 -4453 -2401
rect -4395 -2435 -4379 -2401
rect -4311 -2435 -4295 -2401
rect -4237 -2435 -4221 -2401
rect -4153 -2435 -4137 -2401
rect -4079 -2435 -4063 -2401
rect -3995 -2435 -3979 -2401
rect -3921 -2435 -3905 -2401
rect -3837 -2435 -3821 -2401
rect -3763 -2435 -3747 -2401
rect -3679 -2435 -3663 -2401
rect -3605 -2435 -3589 -2401
rect -3521 -2435 -3505 -2401
rect -3447 -2435 -3431 -2401
rect -3363 -2435 -3347 -2401
rect -3289 -2435 -3273 -2401
rect -3205 -2435 -3189 -2401
rect -3131 -2435 -3115 -2401
rect -3047 -2435 -3031 -2401
rect -2973 -2435 -2957 -2401
rect -2889 -2435 -2873 -2401
rect -2815 -2435 -2799 -2401
rect -2731 -2435 -2715 -2401
rect -2657 -2435 -2641 -2401
rect -2573 -2435 -2557 -2401
rect -2499 -2435 -2483 -2401
rect -2415 -2435 -2399 -2401
rect -2341 -2435 -2325 -2401
rect -2257 -2435 -2241 -2401
rect -2183 -2435 -2167 -2401
rect -2099 -2435 -2083 -2401
rect -2025 -2435 -2009 -2401
rect -1941 -2435 -1925 -2401
rect -1867 -2435 -1851 -2401
rect -1783 -2435 -1767 -2401
rect -1709 -2435 -1693 -2401
rect -1625 -2435 -1609 -2401
rect -1551 -2435 -1535 -2401
rect -1467 -2435 -1451 -2401
rect -1393 -2435 -1377 -2401
rect -1309 -2435 -1293 -2401
rect -1235 -2435 -1219 -2401
rect -1151 -2435 -1135 -2401
rect -1077 -2435 -1061 -2401
rect -993 -2435 -977 -2401
rect -919 -2435 -903 -2401
rect -835 -2435 -819 -2401
rect -761 -2435 -745 -2401
rect -677 -2435 -661 -2401
rect -603 -2435 -587 -2401
rect -519 -2435 -503 -2401
rect -445 -2435 -429 -2401
rect -361 -2435 -345 -2401
rect -287 -2435 -271 -2401
rect -203 -2435 -187 -2401
rect -129 -2435 -113 -2401
rect -45 -2435 -29 -2401
rect 29 -2435 45 -2401
rect 113 -2435 129 -2401
rect 187 -2435 203 -2401
rect 271 -2435 287 -2401
rect 345 -2435 361 -2401
rect 429 -2435 445 -2401
rect 503 -2435 519 -2401
rect 587 -2435 603 -2401
rect 661 -2435 677 -2401
rect 745 -2435 761 -2401
rect 819 -2435 835 -2401
rect 903 -2435 919 -2401
rect 977 -2435 993 -2401
rect 1061 -2435 1077 -2401
rect 1135 -2435 1151 -2401
rect 1219 -2435 1235 -2401
rect 1293 -2435 1309 -2401
rect 1377 -2435 1393 -2401
rect 1451 -2435 1467 -2401
rect 1535 -2435 1551 -2401
rect 1609 -2435 1625 -2401
rect 1693 -2435 1709 -2401
rect 1767 -2435 1783 -2401
rect 1851 -2435 1867 -2401
rect 1925 -2435 1941 -2401
rect 2009 -2435 2025 -2401
rect 2083 -2435 2099 -2401
rect 2167 -2435 2183 -2401
rect 2241 -2435 2257 -2401
rect 2325 -2435 2341 -2401
rect 2399 -2435 2415 -2401
rect 2483 -2435 2499 -2401
rect 2557 -2435 2573 -2401
rect 2641 -2435 2657 -2401
rect 2715 -2435 2731 -2401
rect 2799 -2435 2815 -2401
rect 2873 -2435 2889 -2401
rect 2957 -2435 2973 -2401
rect 3031 -2435 3047 -2401
rect 3115 -2435 3131 -2401
rect 3189 -2435 3205 -2401
rect 3273 -2435 3289 -2401
rect 3347 -2435 3363 -2401
rect 3431 -2435 3447 -2401
rect 3505 -2435 3521 -2401
rect 3589 -2435 3605 -2401
rect 3663 -2435 3679 -2401
rect 3747 -2435 3763 -2401
rect 3821 -2435 3837 -2401
rect 3905 -2435 3921 -2401
rect 3979 -2435 3995 -2401
rect 4063 -2435 4079 -2401
rect 4137 -2435 4153 -2401
rect 4221 -2435 4237 -2401
rect 4295 -2435 4311 -2401
rect 4379 -2435 4395 -2401
rect 4453 -2435 4469 -2401
rect 4537 -2435 4553 -2401
rect 4611 -2435 4627 -2401
rect 4695 -2435 4711 -2401
rect 4769 -2435 4785 -2401
rect 4853 -2435 4869 -2401
rect -5049 -2539 -5015 -2477
rect 5015 -2539 5049 -2477
rect -5049 -2573 -4953 -2539
rect 4953 -2573 5049 -2539
<< viali >>
rect -4853 2401 -4785 2435
rect -4695 2401 -4627 2435
rect -4537 2401 -4469 2435
rect -4379 2401 -4311 2435
rect -4221 2401 -4153 2435
rect -4063 2401 -3995 2435
rect -3905 2401 -3837 2435
rect -3747 2401 -3679 2435
rect -3589 2401 -3521 2435
rect -3431 2401 -3363 2435
rect -3273 2401 -3205 2435
rect -3115 2401 -3047 2435
rect -2957 2401 -2889 2435
rect -2799 2401 -2731 2435
rect -2641 2401 -2573 2435
rect -2483 2401 -2415 2435
rect -2325 2401 -2257 2435
rect -2167 2401 -2099 2435
rect -2009 2401 -1941 2435
rect -1851 2401 -1783 2435
rect -1693 2401 -1625 2435
rect -1535 2401 -1467 2435
rect -1377 2401 -1309 2435
rect -1219 2401 -1151 2435
rect -1061 2401 -993 2435
rect -903 2401 -835 2435
rect -745 2401 -677 2435
rect -587 2401 -519 2435
rect -429 2401 -361 2435
rect -271 2401 -203 2435
rect -113 2401 -45 2435
rect 45 2401 113 2435
rect 203 2401 271 2435
rect 361 2401 429 2435
rect 519 2401 587 2435
rect 677 2401 745 2435
rect 835 2401 903 2435
rect 993 2401 1061 2435
rect 1151 2401 1219 2435
rect 1309 2401 1377 2435
rect 1467 2401 1535 2435
rect 1625 2401 1693 2435
rect 1783 2401 1851 2435
rect 1941 2401 2009 2435
rect 2099 2401 2167 2435
rect 2257 2401 2325 2435
rect 2415 2401 2483 2435
rect 2573 2401 2641 2435
rect 2731 2401 2799 2435
rect 2889 2401 2957 2435
rect 3047 2401 3115 2435
rect 3205 2401 3273 2435
rect 3363 2401 3431 2435
rect 3521 2401 3589 2435
rect 3679 2401 3747 2435
rect 3837 2401 3905 2435
rect 3995 2401 4063 2435
rect 4153 2401 4221 2435
rect 4311 2401 4379 2435
rect 4469 2401 4537 2435
rect 4627 2401 4695 2435
rect 4785 2401 4853 2435
rect -4915 1366 -4881 2342
rect -4757 1366 -4723 2342
rect -4599 1366 -4565 2342
rect -4441 1366 -4407 2342
rect -4283 1366 -4249 2342
rect -4125 1366 -4091 2342
rect -3967 1366 -3933 2342
rect -3809 1366 -3775 2342
rect -3651 1366 -3617 2342
rect -3493 1366 -3459 2342
rect -3335 1366 -3301 2342
rect -3177 1366 -3143 2342
rect -3019 1366 -2985 2342
rect -2861 1366 -2827 2342
rect -2703 1366 -2669 2342
rect -2545 1366 -2511 2342
rect -2387 1366 -2353 2342
rect -2229 1366 -2195 2342
rect -2071 1366 -2037 2342
rect -1913 1366 -1879 2342
rect -1755 1366 -1721 2342
rect -1597 1366 -1563 2342
rect -1439 1366 -1405 2342
rect -1281 1366 -1247 2342
rect -1123 1366 -1089 2342
rect -965 1366 -931 2342
rect -807 1366 -773 2342
rect -649 1366 -615 2342
rect -491 1366 -457 2342
rect -333 1366 -299 2342
rect -175 1366 -141 2342
rect -17 1366 17 2342
rect 141 1366 175 2342
rect 299 1366 333 2342
rect 457 1366 491 2342
rect 615 1366 649 2342
rect 773 1366 807 2342
rect 931 1366 965 2342
rect 1089 1366 1123 2342
rect 1247 1366 1281 2342
rect 1405 1366 1439 2342
rect 1563 1366 1597 2342
rect 1721 1366 1755 2342
rect 1879 1366 1913 2342
rect 2037 1366 2071 2342
rect 2195 1366 2229 2342
rect 2353 1366 2387 2342
rect 2511 1366 2545 2342
rect 2669 1366 2703 2342
rect 2827 1366 2861 2342
rect 2985 1366 3019 2342
rect 3143 1366 3177 2342
rect 3301 1366 3335 2342
rect 3459 1366 3493 2342
rect 3617 1366 3651 2342
rect 3775 1366 3809 2342
rect 3933 1366 3967 2342
rect 4091 1366 4125 2342
rect 4249 1366 4283 2342
rect 4407 1366 4441 2342
rect 4565 1366 4599 2342
rect 4723 1366 4757 2342
rect 4881 1366 4915 2342
rect -4853 1273 -4785 1307
rect -4695 1273 -4627 1307
rect -4537 1273 -4469 1307
rect -4379 1273 -4311 1307
rect -4221 1273 -4153 1307
rect -4063 1273 -3995 1307
rect -3905 1273 -3837 1307
rect -3747 1273 -3679 1307
rect -3589 1273 -3521 1307
rect -3431 1273 -3363 1307
rect -3273 1273 -3205 1307
rect -3115 1273 -3047 1307
rect -2957 1273 -2889 1307
rect -2799 1273 -2731 1307
rect -2641 1273 -2573 1307
rect -2483 1273 -2415 1307
rect -2325 1273 -2257 1307
rect -2167 1273 -2099 1307
rect -2009 1273 -1941 1307
rect -1851 1273 -1783 1307
rect -1693 1273 -1625 1307
rect -1535 1273 -1467 1307
rect -1377 1273 -1309 1307
rect -1219 1273 -1151 1307
rect -1061 1273 -993 1307
rect -903 1273 -835 1307
rect -745 1273 -677 1307
rect -587 1273 -519 1307
rect -429 1273 -361 1307
rect -271 1273 -203 1307
rect -113 1273 -45 1307
rect 45 1273 113 1307
rect 203 1273 271 1307
rect 361 1273 429 1307
rect 519 1273 587 1307
rect 677 1273 745 1307
rect 835 1273 903 1307
rect 993 1273 1061 1307
rect 1151 1273 1219 1307
rect 1309 1273 1377 1307
rect 1467 1273 1535 1307
rect 1625 1273 1693 1307
rect 1783 1273 1851 1307
rect 1941 1273 2009 1307
rect 2099 1273 2167 1307
rect 2257 1273 2325 1307
rect 2415 1273 2483 1307
rect 2573 1273 2641 1307
rect 2731 1273 2799 1307
rect 2889 1273 2957 1307
rect 3047 1273 3115 1307
rect 3205 1273 3273 1307
rect 3363 1273 3431 1307
rect 3521 1273 3589 1307
rect 3679 1273 3747 1307
rect 3837 1273 3905 1307
rect 3995 1273 4063 1307
rect 4153 1273 4221 1307
rect 4311 1273 4379 1307
rect 4469 1273 4537 1307
rect 4627 1273 4695 1307
rect 4785 1273 4853 1307
rect -4853 1165 -4785 1199
rect -4695 1165 -4627 1199
rect -4537 1165 -4469 1199
rect -4379 1165 -4311 1199
rect -4221 1165 -4153 1199
rect -4063 1165 -3995 1199
rect -3905 1165 -3837 1199
rect -3747 1165 -3679 1199
rect -3589 1165 -3521 1199
rect -3431 1165 -3363 1199
rect -3273 1165 -3205 1199
rect -3115 1165 -3047 1199
rect -2957 1165 -2889 1199
rect -2799 1165 -2731 1199
rect -2641 1165 -2573 1199
rect -2483 1165 -2415 1199
rect -2325 1165 -2257 1199
rect -2167 1165 -2099 1199
rect -2009 1165 -1941 1199
rect -1851 1165 -1783 1199
rect -1693 1165 -1625 1199
rect -1535 1165 -1467 1199
rect -1377 1165 -1309 1199
rect -1219 1165 -1151 1199
rect -1061 1165 -993 1199
rect -903 1165 -835 1199
rect -745 1165 -677 1199
rect -587 1165 -519 1199
rect -429 1165 -361 1199
rect -271 1165 -203 1199
rect -113 1165 -45 1199
rect 45 1165 113 1199
rect 203 1165 271 1199
rect 361 1165 429 1199
rect 519 1165 587 1199
rect 677 1165 745 1199
rect 835 1165 903 1199
rect 993 1165 1061 1199
rect 1151 1165 1219 1199
rect 1309 1165 1377 1199
rect 1467 1165 1535 1199
rect 1625 1165 1693 1199
rect 1783 1165 1851 1199
rect 1941 1165 2009 1199
rect 2099 1165 2167 1199
rect 2257 1165 2325 1199
rect 2415 1165 2483 1199
rect 2573 1165 2641 1199
rect 2731 1165 2799 1199
rect 2889 1165 2957 1199
rect 3047 1165 3115 1199
rect 3205 1165 3273 1199
rect 3363 1165 3431 1199
rect 3521 1165 3589 1199
rect 3679 1165 3747 1199
rect 3837 1165 3905 1199
rect 3995 1165 4063 1199
rect 4153 1165 4221 1199
rect 4311 1165 4379 1199
rect 4469 1165 4537 1199
rect 4627 1165 4695 1199
rect 4785 1165 4853 1199
rect -4915 130 -4881 1106
rect -4757 130 -4723 1106
rect -4599 130 -4565 1106
rect -4441 130 -4407 1106
rect -4283 130 -4249 1106
rect -4125 130 -4091 1106
rect -3967 130 -3933 1106
rect -3809 130 -3775 1106
rect -3651 130 -3617 1106
rect -3493 130 -3459 1106
rect -3335 130 -3301 1106
rect -3177 130 -3143 1106
rect -3019 130 -2985 1106
rect -2861 130 -2827 1106
rect -2703 130 -2669 1106
rect -2545 130 -2511 1106
rect -2387 130 -2353 1106
rect -2229 130 -2195 1106
rect -2071 130 -2037 1106
rect -1913 130 -1879 1106
rect -1755 130 -1721 1106
rect -1597 130 -1563 1106
rect -1439 130 -1405 1106
rect -1281 130 -1247 1106
rect -1123 130 -1089 1106
rect -965 130 -931 1106
rect -807 130 -773 1106
rect -649 130 -615 1106
rect -491 130 -457 1106
rect -333 130 -299 1106
rect -175 130 -141 1106
rect -17 130 17 1106
rect 141 130 175 1106
rect 299 130 333 1106
rect 457 130 491 1106
rect 615 130 649 1106
rect 773 130 807 1106
rect 931 130 965 1106
rect 1089 130 1123 1106
rect 1247 130 1281 1106
rect 1405 130 1439 1106
rect 1563 130 1597 1106
rect 1721 130 1755 1106
rect 1879 130 1913 1106
rect 2037 130 2071 1106
rect 2195 130 2229 1106
rect 2353 130 2387 1106
rect 2511 130 2545 1106
rect 2669 130 2703 1106
rect 2827 130 2861 1106
rect 2985 130 3019 1106
rect 3143 130 3177 1106
rect 3301 130 3335 1106
rect 3459 130 3493 1106
rect 3617 130 3651 1106
rect 3775 130 3809 1106
rect 3933 130 3967 1106
rect 4091 130 4125 1106
rect 4249 130 4283 1106
rect 4407 130 4441 1106
rect 4565 130 4599 1106
rect 4723 130 4757 1106
rect 4881 130 4915 1106
rect -4853 37 -4785 71
rect -4695 37 -4627 71
rect -4537 37 -4469 71
rect -4379 37 -4311 71
rect -4221 37 -4153 71
rect -4063 37 -3995 71
rect -3905 37 -3837 71
rect -3747 37 -3679 71
rect -3589 37 -3521 71
rect -3431 37 -3363 71
rect -3273 37 -3205 71
rect -3115 37 -3047 71
rect -2957 37 -2889 71
rect -2799 37 -2731 71
rect -2641 37 -2573 71
rect -2483 37 -2415 71
rect -2325 37 -2257 71
rect -2167 37 -2099 71
rect -2009 37 -1941 71
rect -1851 37 -1783 71
rect -1693 37 -1625 71
rect -1535 37 -1467 71
rect -1377 37 -1309 71
rect -1219 37 -1151 71
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect 1151 37 1219 71
rect 1309 37 1377 71
rect 1467 37 1535 71
rect 1625 37 1693 71
rect 1783 37 1851 71
rect 1941 37 2009 71
rect 2099 37 2167 71
rect 2257 37 2325 71
rect 2415 37 2483 71
rect 2573 37 2641 71
rect 2731 37 2799 71
rect 2889 37 2957 71
rect 3047 37 3115 71
rect 3205 37 3273 71
rect 3363 37 3431 71
rect 3521 37 3589 71
rect 3679 37 3747 71
rect 3837 37 3905 71
rect 3995 37 4063 71
rect 4153 37 4221 71
rect 4311 37 4379 71
rect 4469 37 4537 71
rect 4627 37 4695 71
rect 4785 37 4853 71
rect -4853 -71 -4785 -37
rect -4695 -71 -4627 -37
rect -4537 -71 -4469 -37
rect -4379 -71 -4311 -37
rect -4221 -71 -4153 -37
rect -4063 -71 -3995 -37
rect -3905 -71 -3837 -37
rect -3747 -71 -3679 -37
rect -3589 -71 -3521 -37
rect -3431 -71 -3363 -37
rect -3273 -71 -3205 -37
rect -3115 -71 -3047 -37
rect -2957 -71 -2889 -37
rect -2799 -71 -2731 -37
rect -2641 -71 -2573 -37
rect -2483 -71 -2415 -37
rect -2325 -71 -2257 -37
rect -2167 -71 -2099 -37
rect -2009 -71 -1941 -37
rect -1851 -71 -1783 -37
rect -1693 -71 -1625 -37
rect -1535 -71 -1467 -37
rect -1377 -71 -1309 -37
rect -1219 -71 -1151 -37
rect -1061 -71 -993 -37
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect 993 -71 1061 -37
rect 1151 -71 1219 -37
rect 1309 -71 1377 -37
rect 1467 -71 1535 -37
rect 1625 -71 1693 -37
rect 1783 -71 1851 -37
rect 1941 -71 2009 -37
rect 2099 -71 2167 -37
rect 2257 -71 2325 -37
rect 2415 -71 2483 -37
rect 2573 -71 2641 -37
rect 2731 -71 2799 -37
rect 2889 -71 2957 -37
rect 3047 -71 3115 -37
rect 3205 -71 3273 -37
rect 3363 -71 3431 -37
rect 3521 -71 3589 -37
rect 3679 -71 3747 -37
rect 3837 -71 3905 -37
rect 3995 -71 4063 -37
rect 4153 -71 4221 -37
rect 4311 -71 4379 -37
rect 4469 -71 4537 -37
rect 4627 -71 4695 -37
rect 4785 -71 4853 -37
rect -4915 -1106 -4881 -130
rect -4757 -1106 -4723 -130
rect -4599 -1106 -4565 -130
rect -4441 -1106 -4407 -130
rect -4283 -1106 -4249 -130
rect -4125 -1106 -4091 -130
rect -3967 -1106 -3933 -130
rect -3809 -1106 -3775 -130
rect -3651 -1106 -3617 -130
rect -3493 -1106 -3459 -130
rect -3335 -1106 -3301 -130
rect -3177 -1106 -3143 -130
rect -3019 -1106 -2985 -130
rect -2861 -1106 -2827 -130
rect -2703 -1106 -2669 -130
rect -2545 -1106 -2511 -130
rect -2387 -1106 -2353 -130
rect -2229 -1106 -2195 -130
rect -2071 -1106 -2037 -130
rect -1913 -1106 -1879 -130
rect -1755 -1106 -1721 -130
rect -1597 -1106 -1563 -130
rect -1439 -1106 -1405 -130
rect -1281 -1106 -1247 -130
rect -1123 -1106 -1089 -130
rect -965 -1106 -931 -130
rect -807 -1106 -773 -130
rect -649 -1106 -615 -130
rect -491 -1106 -457 -130
rect -333 -1106 -299 -130
rect -175 -1106 -141 -130
rect -17 -1106 17 -130
rect 141 -1106 175 -130
rect 299 -1106 333 -130
rect 457 -1106 491 -130
rect 615 -1106 649 -130
rect 773 -1106 807 -130
rect 931 -1106 965 -130
rect 1089 -1106 1123 -130
rect 1247 -1106 1281 -130
rect 1405 -1106 1439 -130
rect 1563 -1106 1597 -130
rect 1721 -1106 1755 -130
rect 1879 -1106 1913 -130
rect 2037 -1106 2071 -130
rect 2195 -1106 2229 -130
rect 2353 -1106 2387 -130
rect 2511 -1106 2545 -130
rect 2669 -1106 2703 -130
rect 2827 -1106 2861 -130
rect 2985 -1106 3019 -130
rect 3143 -1106 3177 -130
rect 3301 -1106 3335 -130
rect 3459 -1106 3493 -130
rect 3617 -1106 3651 -130
rect 3775 -1106 3809 -130
rect 3933 -1106 3967 -130
rect 4091 -1106 4125 -130
rect 4249 -1106 4283 -130
rect 4407 -1106 4441 -130
rect 4565 -1106 4599 -130
rect 4723 -1106 4757 -130
rect 4881 -1106 4915 -130
rect -4853 -1199 -4785 -1165
rect -4695 -1199 -4627 -1165
rect -4537 -1199 -4469 -1165
rect -4379 -1199 -4311 -1165
rect -4221 -1199 -4153 -1165
rect -4063 -1199 -3995 -1165
rect -3905 -1199 -3837 -1165
rect -3747 -1199 -3679 -1165
rect -3589 -1199 -3521 -1165
rect -3431 -1199 -3363 -1165
rect -3273 -1199 -3205 -1165
rect -3115 -1199 -3047 -1165
rect -2957 -1199 -2889 -1165
rect -2799 -1199 -2731 -1165
rect -2641 -1199 -2573 -1165
rect -2483 -1199 -2415 -1165
rect -2325 -1199 -2257 -1165
rect -2167 -1199 -2099 -1165
rect -2009 -1199 -1941 -1165
rect -1851 -1199 -1783 -1165
rect -1693 -1199 -1625 -1165
rect -1535 -1199 -1467 -1165
rect -1377 -1199 -1309 -1165
rect -1219 -1199 -1151 -1165
rect -1061 -1199 -993 -1165
rect -903 -1199 -835 -1165
rect -745 -1199 -677 -1165
rect -587 -1199 -519 -1165
rect -429 -1199 -361 -1165
rect -271 -1199 -203 -1165
rect -113 -1199 -45 -1165
rect 45 -1199 113 -1165
rect 203 -1199 271 -1165
rect 361 -1199 429 -1165
rect 519 -1199 587 -1165
rect 677 -1199 745 -1165
rect 835 -1199 903 -1165
rect 993 -1199 1061 -1165
rect 1151 -1199 1219 -1165
rect 1309 -1199 1377 -1165
rect 1467 -1199 1535 -1165
rect 1625 -1199 1693 -1165
rect 1783 -1199 1851 -1165
rect 1941 -1199 2009 -1165
rect 2099 -1199 2167 -1165
rect 2257 -1199 2325 -1165
rect 2415 -1199 2483 -1165
rect 2573 -1199 2641 -1165
rect 2731 -1199 2799 -1165
rect 2889 -1199 2957 -1165
rect 3047 -1199 3115 -1165
rect 3205 -1199 3273 -1165
rect 3363 -1199 3431 -1165
rect 3521 -1199 3589 -1165
rect 3679 -1199 3747 -1165
rect 3837 -1199 3905 -1165
rect 3995 -1199 4063 -1165
rect 4153 -1199 4221 -1165
rect 4311 -1199 4379 -1165
rect 4469 -1199 4537 -1165
rect 4627 -1199 4695 -1165
rect 4785 -1199 4853 -1165
rect -4853 -1307 -4785 -1273
rect -4695 -1307 -4627 -1273
rect -4537 -1307 -4469 -1273
rect -4379 -1307 -4311 -1273
rect -4221 -1307 -4153 -1273
rect -4063 -1307 -3995 -1273
rect -3905 -1307 -3837 -1273
rect -3747 -1307 -3679 -1273
rect -3589 -1307 -3521 -1273
rect -3431 -1307 -3363 -1273
rect -3273 -1307 -3205 -1273
rect -3115 -1307 -3047 -1273
rect -2957 -1307 -2889 -1273
rect -2799 -1307 -2731 -1273
rect -2641 -1307 -2573 -1273
rect -2483 -1307 -2415 -1273
rect -2325 -1307 -2257 -1273
rect -2167 -1307 -2099 -1273
rect -2009 -1307 -1941 -1273
rect -1851 -1307 -1783 -1273
rect -1693 -1307 -1625 -1273
rect -1535 -1307 -1467 -1273
rect -1377 -1307 -1309 -1273
rect -1219 -1307 -1151 -1273
rect -1061 -1307 -993 -1273
rect -903 -1307 -835 -1273
rect -745 -1307 -677 -1273
rect -587 -1307 -519 -1273
rect -429 -1307 -361 -1273
rect -271 -1307 -203 -1273
rect -113 -1307 -45 -1273
rect 45 -1307 113 -1273
rect 203 -1307 271 -1273
rect 361 -1307 429 -1273
rect 519 -1307 587 -1273
rect 677 -1307 745 -1273
rect 835 -1307 903 -1273
rect 993 -1307 1061 -1273
rect 1151 -1307 1219 -1273
rect 1309 -1307 1377 -1273
rect 1467 -1307 1535 -1273
rect 1625 -1307 1693 -1273
rect 1783 -1307 1851 -1273
rect 1941 -1307 2009 -1273
rect 2099 -1307 2167 -1273
rect 2257 -1307 2325 -1273
rect 2415 -1307 2483 -1273
rect 2573 -1307 2641 -1273
rect 2731 -1307 2799 -1273
rect 2889 -1307 2957 -1273
rect 3047 -1307 3115 -1273
rect 3205 -1307 3273 -1273
rect 3363 -1307 3431 -1273
rect 3521 -1307 3589 -1273
rect 3679 -1307 3747 -1273
rect 3837 -1307 3905 -1273
rect 3995 -1307 4063 -1273
rect 4153 -1307 4221 -1273
rect 4311 -1307 4379 -1273
rect 4469 -1307 4537 -1273
rect 4627 -1307 4695 -1273
rect 4785 -1307 4853 -1273
rect -4915 -2342 -4881 -1366
rect -4757 -2342 -4723 -1366
rect -4599 -2342 -4565 -1366
rect -4441 -2342 -4407 -1366
rect -4283 -2342 -4249 -1366
rect -4125 -2342 -4091 -1366
rect -3967 -2342 -3933 -1366
rect -3809 -2342 -3775 -1366
rect -3651 -2342 -3617 -1366
rect -3493 -2342 -3459 -1366
rect -3335 -2342 -3301 -1366
rect -3177 -2342 -3143 -1366
rect -3019 -2342 -2985 -1366
rect -2861 -2342 -2827 -1366
rect -2703 -2342 -2669 -1366
rect -2545 -2342 -2511 -1366
rect -2387 -2342 -2353 -1366
rect -2229 -2342 -2195 -1366
rect -2071 -2342 -2037 -1366
rect -1913 -2342 -1879 -1366
rect -1755 -2342 -1721 -1366
rect -1597 -2342 -1563 -1366
rect -1439 -2342 -1405 -1366
rect -1281 -2342 -1247 -1366
rect -1123 -2342 -1089 -1366
rect -965 -2342 -931 -1366
rect -807 -2342 -773 -1366
rect -649 -2342 -615 -1366
rect -491 -2342 -457 -1366
rect -333 -2342 -299 -1366
rect -175 -2342 -141 -1366
rect -17 -2342 17 -1366
rect 141 -2342 175 -1366
rect 299 -2342 333 -1366
rect 457 -2342 491 -1366
rect 615 -2342 649 -1366
rect 773 -2342 807 -1366
rect 931 -2342 965 -1366
rect 1089 -2342 1123 -1366
rect 1247 -2342 1281 -1366
rect 1405 -2342 1439 -1366
rect 1563 -2342 1597 -1366
rect 1721 -2342 1755 -1366
rect 1879 -2342 1913 -1366
rect 2037 -2342 2071 -1366
rect 2195 -2342 2229 -1366
rect 2353 -2342 2387 -1366
rect 2511 -2342 2545 -1366
rect 2669 -2342 2703 -1366
rect 2827 -2342 2861 -1366
rect 2985 -2342 3019 -1366
rect 3143 -2342 3177 -1366
rect 3301 -2342 3335 -1366
rect 3459 -2342 3493 -1366
rect 3617 -2342 3651 -1366
rect 3775 -2342 3809 -1366
rect 3933 -2342 3967 -1366
rect 4091 -2342 4125 -1366
rect 4249 -2342 4283 -1366
rect 4407 -2342 4441 -1366
rect 4565 -2342 4599 -1366
rect 4723 -2342 4757 -1366
rect 4881 -2342 4915 -1366
rect -4853 -2435 -4785 -2401
rect -4695 -2435 -4627 -2401
rect -4537 -2435 -4469 -2401
rect -4379 -2435 -4311 -2401
rect -4221 -2435 -4153 -2401
rect -4063 -2435 -3995 -2401
rect -3905 -2435 -3837 -2401
rect -3747 -2435 -3679 -2401
rect -3589 -2435 -3521 -2401
rect -3431 -2435 -3363 -2401
rect -3273 -2435 -3205 -2401
rect -3115 -2435 -3047 -2401
rect -2957 -2435 -2889 -2401
rect -2799 -2435 -2731 -2401
rect -2641 -2435 -2573 -2401
rect -2483 -2435 -2415 -2401
rect -2325 -2435 -2257 -2401
rect -2167 -2435 -2099 -2401
rect -2009 -2435 -1941 -2401
rect -1851 -2435 -1783 -2401
rect -1693 -2435 -1625 -2401
rect -1535 -2435 -1467 -2401
rect -1377 -2435 -1309 -2401
rect -1219 -2435 -1151 -2401
rect -1061 -2435 -993 -2401
rect -903 -2435 -835 -2401
rect -745 -2435 -677 -2401
rect -587 -2435 -519 -2401
rect -429 -2435 -361 -2401
rect -271 -2435 -203 -2401
rect -113 -2435 -45 -2401
rect 45 -2435 113 -2401
rect 203 -2435 271 -2401
rect 361 -2435 429 -2401
rect 519 -2435 587 -2401
rect 677 -2435 745 -2401
rect 835 -2435 903 -2401
rect 993 -2435 1061 -2401
rect 1151 -2435 1219 -2401
rect 1309 -2435 1377 -2401
rect 1467 -2435 1535 -2401
rect 1625 -2435 1693 -2401
rect 1783 -2435 1851 -2401
rect 1941 -2435 2009 -2401
rect 2099 -2435 2167 -2401
rect 2257 -2435 2325 -2401
rect 2415 -2435 2483 -2401
rect 2573 -2435 2641 -2401
rect 2731 -2435 2799 -2401
rect 2889 -2435 2957 -2401
rect 3047 -2435 3115 -2401
rect 3205 -2435 3273 -2401
rect 3363 -2435 3431 -2401
rect 3521 -2435 3589 -2401
rect 3679 -2435 3747 -2401
rect 3837 -2435 3905 -2401
rect 3995 -2435 4063 -2401
rect 4153 -2435 4221 -2401
rect 4311 -2435 4379 -2401
rect 4469 -2435 4537 -2401
rect 4627 -2435 4695 -2401
rect 4785 -2435 4853 -2401
<< metal1 >>
rect -4865 2435 -4773 2441
rect -4865 2401 -4853 2435
rect -4785 2401 -4773 2435
rect -4865 2395 -4773 2401
rect -4707 2435 -4615 2441
rect -4707 2401 -4695 2435
rect -4627 2401 -4615 2435
rect -4707 2395 -4615 2401
rect -4549 2435 -4457 2441
rect -4549 2401 -4537 2435
rect -4469 2401 -4457 2435
rect -4549 2395 -4457 2401
rect -4391 2435 -4299 2441
rect -4391 2401 -4379 2435
rect -4311 2401 -4299 2435
rect -4391 2395 -4299 2401
rect -4233 2435 -4141 2441
rect -4233 2401 -4221 2435
rect -4153 2401 -4141 2435
rect -4233 2395 -4141 2401
rect -4075 2435 -3983 2441
rect -4075 2401 -4063 2435
rect -3995 2401 -3983 2435
rect -4075 2395 -3983 2401
rect -3917 2435 -3825 2441
rect -3917 2401 -3905 2435
rect -3837 2401 -3825 2435
rect -3917 2395 -3825 2401
rect -3759 2435 -3667 2441
rect -3759 2401 -3747 2435
rect -3679 2401 -3667 2435
rect -3759 2395 -3667 2401
rect -3601 2435 -3509 2441
rect -3601 2401 -3589 2435
rect -3521 2401 -3509 2435
rect -3601 2395 -3509 2401
rect -3443 2435 -3351 2441
rect -3443 2401 -3431 2435
rect -3363 2401 -3351 2435
rect -3443 2395 -3351 2401
rect -3285 2435 -3193 2441
rect -3285 2401 -3273 2435
rect -3205 2401 -3193 2435
rect -3285 2395 -3193 2401
rect -3127 2435 -3035 2441
rect -3127 2401 -3115 2435
rect -3047 2401 -3035 2435
rect -3127 2395 -3035 2401
rect -2969 2435 -2877 2441
rect -2969 2401 -2957 2435
rect -2889 2401 -2877 2435
rect -2969 2395 -2877 2401
rect -2811 2435 -2719 2441
rect -2811 2401 -2799 2435
rect -2731 2401 -2719 2435
rect -2811 2395 -2719 2401
rect -2653 2435 -2561 2441
rect -2653 2401 -2641 2435
rect -2573 2401 -2561 2435
rect -2653 2395 -2561 2401
rect -2495 2435 -2403 2441
rect -2495 2401 -2483 2435
rect -2415 2401 -2403 2435
rect -2495 2395 -2403 2401
rect -2337 2435 -2245 2441
rect -2337 2401 -2325 2435
rect -2257 2401 -2245 2435
rect -2337 2395 -2245 2401
rect -2179 2435 -2087 2441
rect -2179 2401 -2167 2435
rect -2099 2401 -2087 2435
rect -2179 2395 -2087 2401
rect -2021 2435 -1929 2441
rect -2021 2401 -2009 2435
rect -1941 2401 -1929 2435
rect -2021 2395 -1929 2401
rect -1863 2435 -1771 2441
rect -1863 2401 -1851 2435
rect -1783 2401 -1771 2435
rect -1863 2395 -1771 2401
rect -1705 2435 -1613 2441
rect -1705 2401 -1693 2435
rect -1625 2401 -1613 2435
rect -1705 2395 -1613 2401
rect -1547 2435 -1455 2441
rect -1547 2401 -1535 2435
rect -1467 2401 -1455 2435
rect -1547 2395 -1455 2401
rect -1389 2435 -1297 2441
rect -1389 2401 -1377 2435
rect -1309 2401 -1297 2435
rect -1389 2395 -1297 2401
rect -1231 2435 -1139 2441
rect -1231 2401 -1219 2435
rect -1151 2401 -1139 2435
rect -1231 2395 -1139 2401
rect -1073 2435 -981 2441
rect -1073 2401 -1061 2435
rect -993 2401 -981 2435
rect -1073 2395 -981 2401
rect -915 2435 -823 2441
rect -915 2401 -903 2435
rect -835 2401 -823 2435
rect -915 2395 -823 2401
rect -757 2435 -665 2441
rect -757 2401 -745 2435
rect -677 2401 -665 2435
rect -757 2395 -665 2401
rect -599 2435 -507 2441
rect -599 2401 -587 2435
rect -519 2401 -507 2435
rect -599 2395 -507 2401
rect -441 2435 -349 2441
rect -441 2401 -429 2435
rect -361 2401 -349 2435
rect -441 2395 -349 2401
rect -283 2435 -191 2441
rect -283 2401 -271 2435
rect -203 2401 -191 2435
rect -283 2395 -191 2401
rect -125 2435 -33 2441
rect -125 2401 -113 2435
rect -45 2401 -33 2435
rect -125 2395 -33 2401
rect 33 2435 125 2441
rect 33 2401 45 2435
rect 113 2401 125 2435
rect 33 2395 125 2401
rect 191 2435 283 2441
rect 191 2401 203 2435
rect 271 2401 283 2435
rect 191 2395 283 2401
rect 349 2435 441 2441
rect 349 2401 361 2435
rect 429 2401 441 2435
rect 349 2395 441 2401
rect 507 2435 599 2441
rect 507 2401 519 2435
rect 587 2401 599 2435
rect 507 2395 599 2401
rect 665 2435 757 2441
rect 665 2401 677 2435
rect 745 2401 757 2435
rect 665 2395 757 2401
rect 823 2435 915 2441
rect 823 2401 835 2435
rect 903 2401 915 2435
rect 823 2395 915 2401
rect 981 2435 1073 2441
rect 981 2401 993 2435
rect 1061 2401 1073 2435
rect 981 2395 1073 2401
rect 1139 2435 1231 2441
rect 1139 2401 1151 2435
rect 1219 2401 1231 2435
rect 1139 2395 1231 2401
rect 1297 2435 1389 2441
rect 1297 2401 1309 2435
rect 1377 2401 1389 2435
rect 1297 2395 1389 2401
rect 1455 2435 1547 2441
rect 1455 2401 1467 2435
rect 1535 2401 1547 2435
rect 1455 2395 1547 2401
rect 1613 2435 1705 2441
rect 1613 2401 1625 2435
rect 1693 2401 1705 2435
rect 1613 2395 1705 2401
rect 1771 2435 1863 2441
rect 1771 2401 1783 2435
rect 1851 2401 1863 2435
rect 1771 2395 1863 2401
rect 1929 2435 2021 2441
rect 1929 2401 1941 2435
rect 2009 2401 2021 2435
rect 1929 2395 2021 2401
rect 2087 2435 2179 2441
rect 2087 2401 2099 2435
rect 2167 2401 2179 2435
rect 2087 2395 2179 2401
rect 2245 2435 2337 2441
rect 2245 2401 2257 2435
rect 2325 2401 2337 2435
rect 2245 2395 2337 2401
rect 2403 2435 2495 2441
rect 2403 2401 2415 2435
rect 2483 2401 2495 2435
rect 2403 2395 2495 2401
rect 2561 2435 2653 2441
rect 2561 2401 2573 2435
rect 2641 2401 2653 2435
rect 2561 2395 2653 2401
rect 2719 2435 2811 2441
rect 2719 2401 2731 2435
rect 2799 2401 2811 2435
rect 2719 2395 2811 2401
rect 2877 2435 2969 2441
rect 2877 2401 2889 2435
rect 2957 2401 2969 2435
rect 2877 2395 2969 2401
rect 3035 2435 3127 2441
rect 3035 2401 3047 2435
rect 3115 2401 3127 2435
rect 3035 2395 3127 2401
rect 3193 2435 3285 2441
rect 3193 2401 3205 2435
rect 3273 2401 3285 2435
rect 3193 2395 3285 2401
rect 3351 2435 3443 2441
rect 3351 2401 3363 2435
rect 3431 2401 3443 2435
rect 3351 2395 3443 2401
rect 3509 2435 3601 2441
rect 3509 2401 3521 2435
rect 3589 2401 3601 2435
rect 3509 2395 3601 2401
rect 3667 2435 3759 2441
rect 3667 2401 3679 2435
rect 3747 2401 3759 2435
rect 3667 2395 3759 2401
rect 3825 2435 3917 2441
rect 3825 2401 3837 2435
rect 3905 2401 3917 2435
rect 3825 2395 3917 2401
rect 3983 2435 4075 2441
rect 3983 2401 3995 2435
rect 4063 2401 4075 2435
rect 3983 2395 4075 2401
rect 4141 2435 4233 2441
rect 4141 2401 4153 2435
rect 4221 2401 4233 2435
rect 4141 2395 4233 2401
rect 4299 2435 4391 2441
rect 4299 2401 4311 2435
rect 4379 2401 4391 2435
rect 4299 2395 4391 2401
rect 4457 2435 4549 2441
rect 4457 2401 4469 2435
rect 4537 2401 4549 2435
rect 4457 2395 4549 2401
rect 4615 2435 4707 2441
rect 4615 2401 4627 2435
rect 4695 2401 4707 2435
rect 4615 2395 4707 2401
rect 4773 2435 4865 2441
rect 4773 2401 4785 2435
rect 4853 2401 4865 2435
rect 4773 2395 4865 2401
rect -4921 2342 -4875 2354
rect -4921 1366 -4915 2342
rect -4881 1366 -4875 2342
rect -4921 1354 -4875 1366
rect -4763 2342 -4717 2354
rect -4763 1366 -4757 2342
rect -4723 1366 -4717 2342
rect -4763 1354 -4717 1366
rect -4605 2342 -4559 2354
rect -4605 1366 -4599 2342
rect -4565 1366 -4559 2342
rect -4605 1354 -4559 1366
rect -4447 2342 -4401 2354
rect -4447 1366 -4441 2342
rect -4407 1366 -4401 2342
rect -4447 1354 -4401 1366
rect -4289 2342 -4243 2354
rect -4289 1366 -4283 2342
rect -4249 1366 -4243 2342
rect -4289 1354 -4243 1366
rect -4131 2342 -4085 2354
rect -4131 1366 -4125 2342
rect -4091 1366 -4085 2342
rect -4131 1354 -4085 1366
rect -3973 2342 -3927 2354
rect -3973 1366 -3967 2342
rect -3933 1366 -3927 2342
rect -3973 1354 -3927 1366
rect -3815 2342 -3769 2354
rect -3815 1366 -3809 2342
rect -3775 1366 -3769 2342
rect -3815 1354 -3769 1366
rect -3657 2342 -3611 2354
rect -3657 1366 -3651 2342
rect -3617 1366 -3611 2342
rect -3657 1354 -3611 1366
rect -3499 2342 -3453 2354
rect -3499 1366 -3493 2342
rect -3459 1366 -3453 2342
rect -3499 1354 -3453 1366
rect -3341 2342 -3295 2354
rect -3341 1366 -3335 2342
rect -3301 1366 -3295 2342
rect -3341 1354 -3295 1366
rect -3183 2342 -3137 2354
rect -3183 1366 -3177 2342
rect -3143 1366 -3137 2342
rect -3183 1354 -3137 1366
rect -3025 2342 -2979 2354
rect -3025 1366 -3019 2342
rect -2985 1366 -2979 2342
rect -3025 1354 -2979 1366
rect -2867 2342 -2821 2354
rect -2867 1366 -2861 2342
rect -2827 1366 -2821 2342
rect -2867 1354 -2821 1366
rect -2709 2342 -2663 2354
rect -2709 1366 -2703 2342
rect -2669 1366 -2663 2342
rect -2709 1354 -2663 1366
rect -2551 2342 -2505 2354
rect -2551 1366 -2545 2342
rect -2511 1366 -2505 2342
rect -2551 1354 -2505 1366
rect -2393 2342 -2347 2354
rect -2393 1366 -2387 2342
rect -2353 1366 -2347 2342
rect -2393 1354 -2347 1366
rect -2235 2342 -2189 2354
rect -2235 1366 -2229 2342
rect -2195 1366 -2189 2342
rect -2235 1354 -2189 1366
rect -2077 2342 -2031 2354
rect -2077 1366 -2071 2342
rect -2037 1366 -2031 2342
rect -2077 1354 -2031 1366
rect -1919 2342 -1873 2354
rect -1919 1366 -1913 2342
rect -1879 1366 -1873 2342
rect -1919 1354 -1873 1366
rect -1761 2342 -1715 2354
rect -1761 1366 -1755 2342
rect -1721 1366 -1715 2342
rect -1761 1354 -1715 1366
rect -1603 2342 -1557 2354
rect -1603 1366 -1597 2342
rect -1563 1366 -1557 2342
rect -1603 1354 -1557 1366
rect -1445 2342 -1399 2354
rect -1445 1366 -1439 2342
rect -1405 1366 -1399 2342
rect -1445 1354 -1399 1366
rect -1287 2342 -1241 2354
rect -1287 1366 -1281 2342
rect -1247 1366 -1241 2342
rect -1287 1354 -1241 1366
rect -1129 2342 -1083 2354
rect -1129 1366 -1123 2342
rect -1089 1366 -1083 2342
rect -1129 1354 -1083 1366
rect -971 2342 -925 2354
rect -971 1366 -965 2342
rect -931 1366 -925 2342
rect -971 1354 -925 1366
rect -813 2342 -767 2354
rect -813 1366 -807 2342
rect -773 1366 -767 2342
rect -813 1354 -767 1366
rect -655 2342 -609 2354
rect -655 1366 -649 2342
rect -615 1366 -609 2342
rect -655 1354 -609 1366
rect -497 2342 -451 2354
rect -497 1366 -491 2342
rect -457 1366 -451 2342
rect -497 1354 -451 1366
rect -339 2342 -293 2354
rect -339 1366 -333 2342
rect -299 1366 -293 2342
rect -339 1354 -293 1366
rect -181 2342 -135 2354
rect -181 1366 -175 2342
rect -141 1366 -135 2342
rect -181 1354 -135 1366
rect -23 2342 23 2354
rect -23 1366 -17 2342
rect 17 1366 23 2342
rect -23 1354 23 1366
rect 135 2342 181 2354
rect 135 1366 141 2342
rect 175 1366 181 2342
rect 135 1354 181 1366
rect 293 2342 339 2354
rect 293 1366 299 2342
rect 333 1366 339 2342
rect 293 1354 339 1366
rect 451 2342 497 2354
rect 451 1366 457 2342
rect 491 1366 497 2342
rect 451 1354 497 1366
rect 609 2342 655 2354
rect 609 1366 615 2342
rect 649 1366 655 2342
rect 609 1354 655 1366
rect 767 2342 813 2354
rect 767 1366 773 2342
rect 807 1366 813 2342
rect 767 1354 813 1366
rect 925 2342 971 2354
rect 925 1366 931 2342
rect 965 1366 971 2342
rect 925 1354 971 1366
rect 1083 2342 1129 2354
rect 1083 1366 1089 2342
rect 1123 1366 1129 2342
rect 1083 1354 1129 1366
rect 1241 2342 1287 2354
rect 1241 1366 1247 2342
rect 1281 1366 1287 2342
rect 1241 1354 1287 1366
rect 1399 2342 1445 2354
rect 1399 1366 1405 2342
rect 1439 1366 1445 2342
rect 1399 1354 1445 1366
rect 1557 2342 1603 2354
rect 1557 1366 1563 2342
rect 1597 1366 1603 2342
rect 1557 1354 1603 1366
rect 1715 2342 1761 2354
rect 1715 1366 1721 2342
rect 1755 1366 1761 2342
rect 1715 1354 1761 1366
rect 1873 2342 1919 2354
rect 1873 1366 1879 2342
rect 1913 1366 1919 2342
rect 1873 1354 1919 1366
rect 2031 2342 2077 2354
rect 2031 1366 2037 2342
rect 2071 1366 2077 2342
rect 2031 1354 2077 1366
rect 2189 2342 2235 2354
rect 2189 1366 2195 2342
rect 2229 1366 2235 2342
rect 2189 1354 2235 1366
rect 2347 2342 2393 2354
rect 2347 1366 2353 2342
rect 2387 1366 2393 2342
rect 2347 1354 2393 1366
rect 2505 2342 2551 2354
rect 2505 1366 2511 2342
rect 2545 1366 2551 2342
rect 2505 1354 2551 1366
rect 2663 2342 2709 2354
rect 2663 1366 2669 2342
rect 2703 1366 2709 2342
rect 2663 1354 2709 1366
rect 2821 2342 2867 2354
rect 2821 1366 2827 2342
rect 2861 1366 2867 2342
rect 2821 1354 2867 1366
rect 2979 2342 3025 2354
rect 2979 1366 2985 2342
rect 3019 1366 3025 2342
rect 2979 1354 3025 1366
rect 3137 2342 3183 2354
rect 3137 1366 3143 2342
rect 3177 1366 3183 2342
rect 3137 1354 3183 1366
rect 3295 2342 3341 2354
rect 3295 1366 3301 2342
rect 3335 1366 3341 2342
rect 3295 1354 3341 1366
rect 3453 2342 3499 2354
rect 3453 1366 3459 2342
rect 3493 1366 3499 2342
rect 3453 1354 3499 1366
rect 3611 2342 3657 2354
rect 3611 1366 3617 2342
rect 3651 1366 3657 2342
rect 3611 1354 3657 1366
rect 3769 2342 3815 2354
rect 3769 1366 3775 2342
rect 3809 1366 3815 2342
rect 3769 1354 3815 1366
rect 3927 2342 3973 2354
rect 3927 1366 3933 2342
rect 3967 1366 3973 2342
rect 3927 1354 3973 1366
rect 4085 2342 4131 2354
rect 4085 1366 4091 2342
rect 4125 1366 4131 2342
rect 4085 1354 4131 1366
rect 4243 2342 4289 2354
rect 4243 1366 4249 2342
rect 4283 1366 4289 2342
rect 4243 1354 4289 1366
rect 4401 2342 4447 2354
rect 4401 1366 4407 2342
rect 4441 1366 4447 2342
rect 4401 1354 4447 1366
rect 4559 2342 4605 2354
rect 4559 1366 4565 2342
rect 4599 1366 4605 2342
rect 4559 1354 4605 1366
rect 4717 2342 4763 2354
rect 4717 1366 4723 2342
rect 4757 1366 4763 2342
rect 4717 1354 4763 1366
rect 4875 2342 4921 2354
rect 4875 1366 4881 2342
rect 4915 1366 4921 2342
rect 4875 1354 4921 1366
rect -4865 1307 -4773 1313
rect -4865 1273 -4853 1307
rect -4785 1273 -4773 1307
rect -4865 1267 -4773 1273
rect -4707 1307 -4615 1313
rect -4707 1273 -4695 1307
rect -4627 1273 -4615 1307
rect -4707 1267 -4615 1273
rect -4549 1307 -4457 1313
rect -4549 1273 -4537 1307
rect -4469 1273 -4457 1307
rect -4549 1267 -4457 1273
rect -4391 1307 -4299 1313
rect -4391 1273 -4379 1307
rect -4311 1273 -4299 1307
rect -4391 1267 -4299 1273
rect -4233 1307 -4141 1313
rect -4233 1273 -4221 1307
rect -4153 1273 -4141 1307
rect -4233 1267 -4141 1273
rect -4075 1307 -3983 1313
rect -4075 1273 -4063 1307
rect -3995 1273 -3983 1307
rect -4075 1267 -3983 1273
rect -3917 1307 -3825 1313
rect -3917 1273 -3905 1307
rect -3837 1273 -3825 1307
rect -3917 1267 -3825 1273
rect -3759 1307 -3667 1313
rect -3759 1273 -3747 1307
rect -3679 1273 -3667 1307
rect -3759 1267 -3667 1273
rect -3601 1307 -3509 1313
rect -3601 1273 -3589 1307
rect -3521 1273 -3509 1307
rect -3601 1267 -3509 1273
rect -3443 1307 -3351 1313
rect -3443 1273 -3431 1307
rect -3363 1273 -3351 1307
rect -3443 1267 -3351 1273
rect -3285 1307 -3193 1313
rect -3285 1273 -3273 1307
rect -3205 1273 -3193 1307
rect -3285 1267 -3193 1273
rect -3127 1307 -3035 1313
rect -3127 1273 -3115 1307
rect -3047 1273 -3035 1307
rect -3127 1267 -3035 1273
rect -2969 1307 -2877 1313
rect -2969 1273 -2957 1307
rect -2889 1273 -2877 1307
rect -2969 1267 -2877 1273
rect -2811 1307 -2719 1313
rect -2811 1273 -2799 1307
rect -2731 1273 -2719 1307
rect -2811 1267 -2719 1273
rect -2653 1307 -2561 1313
rect -2653 1273 -2641 1307
rect -2573 1273 -2561 1307
rect -2653 1267 -2561 1273
rect -2495 1307 -2403 1313
rect -2495 1273 -2483 1307
rect -2415 1273 -2403 1307
rect -2495 1267 -2403 1273
rect -2337 1307 -2245 1313
rect -2337 1273 -2325 1307
rect -2257 1273 -2245 1307
rect -2337 1267 -2245 1273
rect -2179 1307 -2087 1313
rect -2179 1273 -2167 1307
rect -2099 1273 -2087 1307
rect -2179 1267 -2087 1273
rect -2021 1307 -1929 1313
rect -2021 1273 -2009 1307
rect -1941 1273 -1929 1307
rect -2021 1267 -1929 1273
rect -1863 1307 -1771 1313
rect -1863 1273 -1851 1307
rect -1783 1273 -1771 1307
rect -1863 1267 -1771 1273
rect -1705 1307 -1613 1313
rect -1705 1273 -1693 1307
rect -1625 1273 -1613 1307
rect -1705 1267 -1613 1273
rect -1547 1307 -1455 1313
rect -1547 1273 -1535 1307
rect -1467 1273 -1455 1307
rect -1547 1267 -1455 1273
rect -1389 1307 -1297 1313
rect -1389 1273 -1377 1307
rect -1309 1273 -1297 1307
rect -1389 1267 -1297 1273
rect -1231 1307 -1139 1313
rect -1231 1273 -1219 1307
rect -1151 1273 -1139 1307
rect -1231 1267 -1139 1273
rect -1073 1307 -981 1313
rect -1073 1273 -1061 1307
rect -993 1273 -981 1307
rect -1073 1267 -981 1273
rect -915 1307 -823 1313
rect -915 1273 -903 1307
rect -835 1273 -823 1307
rect -915 1267 -823 1273
rect -757 1307 -665 1313
rect -757 1273 -745 1307
rect -677 1273 -665 1307
rect -757 1267 -665 1273
rect -599 1307 -507 1313
rect -599 1273 -587 1307
rect -519 1273 -507 1307
rect -599 1267 -507 1273
rect -441 1307 -349 1313
rect -441 1273 -429 1307
rect -361 1273 -349 1307
rect -441 1267 -349 1273
rect -283 1307 -191 1313
rect -283 1273 -271 1307
rect -203 1273 -191 1307
rect -283 1267 -191 1273
rect -125 1307 -33 1313
rect -125 1273 -113 1307
rect -45 1273 -33 1307
rect -125 1267 -33 1273
rect 33 1307 125 1313
rect 33 1273 45 1307
rect 113 1273 125 1307
rect 33 1267 125 1273
rect 191 1307 283 1313
rect 191 1273 203 1307
rect 271 1273 283 1307
rect 191 1267 283 1273
rect 349 1307 441 1313
rect 349 1273 361 1307
rect 429 1273 441 1307
rect 349 1267 441 1273
rect 507 1307 599 1313
rect 507 1273 519 1307
rect 587 1273 599 1307
rect 507 1267 599 1273
rect 665 1307 757 1313
rect 665 1273 677 1307
rect 745 1273 757 1307
rect 665 1267 757 1273
rect 823 1307 915 1313
rect 823 1273 835 1307
rect 903 1273 915 1307
rect 823 1267 915 1273
rect 981 1307 1073 1313
rect 981 1273 993 1307
rect 1061 1273 1073 1307
rect 981 1267 1073 1273
rect 1139 1307 1231 1313
rect 1139 1273 1151 1307
rect 1219 1273 1231 1307
rect 1139 1267 1231 1273
rect 1297 1307 1389 1313
rect 1297 1273 1309 1307
rect 1377 1273 1389 1307
rect 1297 1267 1389 1273
rect 1455 1307 1547 1313
rect 1455 1273 1467 1307
rect 1535 1273 1547 1307
rect 1455 1267 1547 1273
rect 1613 1307 1705 1313
rect 1613 1273 1625 1307
rect 1693 1273 1705 1307
rect 1613 1267 1705 1273
rect 1771 1307 1863 1313
rect 1771 1273 1783 1307
rect 1851 1273 1863 1307
rect 1771 1267 1863 1273
rect 1929 1307 2021 1313
rect 1929 1273 1941 1307
rect 2009 1273 2021 1307
rect 1929 1267 2021 1273
rect 2087 1307 2179 1313
rect 2087 1273 2099 1307
rect 2167 1273 2179 1307
rect 2087 1267 2179 1273
rect 2245 1307 2337 1313
rect 2245 1273 2257 1307
rect 2325 1273 2337 1307
rect 2245 1267 2337 1273
rect 2403 1307 2495 1313
rect 2403 1273 2415 1307
rect 2483 1273 2495 1307
rect 2403 1267 2495 1273
rect 2561 1307 2653 1313
rect 2561 1273 2573 1307
rect 2641 1273 2653 1307
rect 2561 1267 2653 1273
rect 2719 1307 2811 1313
rect 2719 1273 2731 1307
rect 2799 1273 2811 1307
rect 2719 1267 2811 1273
rect 2877 1307 2969 1313
rect 2877 1273 2889 1307
rect 2957 1273 2969 1307
rect 2877 1267 2969 1273
rect 3035 1307 3127 1313
rect 3035 1273 3047 1307
rect 3115 1273 3127 1307
rect 3035 1267 3127 1273
rect 3193 1307 3285 1313
rect 3193 1273 3205 1307
rect 3273 1273 3285 1307
rect 3193 1267 3285 1273
rect 3351 1307 3443 1313
rect 3351 1273 3363 1307
rect 3431 1273 3443 1307
rect 3351 1267 3443 1273
rect 3509 1307 3601 1313
rect 3509 1273 3521 1307
rect 3589 1273 3601 1307
rect 3509 1267 3601 1273
rect 3667 1307 3759 1313
rect 3667 1273 3679 1307
rect 3747 1273 3759 1307
rect 3667 1267 3759 1273
rect 3825 1307 3917 1313
rect 3825 1273 3837 1307
rect 3905 1273 3917 1307
rect 3825 1267 3917 1273
rect 3983 1307 4075 1313
rect 3983 1273 3995 1307
rect 4063 1273 4075 1307
rect 3983 1267 4075 1273
rect 4141 1307 4233 1313
rect 4141 1273 4153 1307
rect 4221 1273 4233 1307
rect 4141 1267 4233 1273
rect 4299 1307 4391 1313
rect 4299 1273 4311 1307
rect 4379 1273 4391 1307
rect 4299 1267 4391 1273
rect 4457 1307 4549 1313
rect 4457 1273 4469 1307
rect 4537 1273 4549 1307
rect 4457 1267 4549 1273
rect 4615 1307 4707 1313
rect 4615 1273 4627 1307
rect 4695 1273 4707 1307
rect 4615 1267 4707 1273
rect 4773 1307 4865 1313
rect 4773 1273 4785 1307
rect 4853 1273 4865 1307
rect 4773 1267 4865 1273
rect -4865 1199 -4773 1205
rect -4865 1165 -4853 1199
rect -4785 1165 -4773 1199
rect -4865 1159 -4773 1165
rect -4707 1199 -4615 1205
rect -4707 1165 -4695 1199
rect -4627 1165 -4615 1199
rect -4707 1159 -4615 1165
rect -4549 1199 -4457 1205
rect -4549 1165 -4537 1199
rect -4469 1165 -4457 1199
rect -4549 1159 -4457 1165
rect -4391 1199 -4299 1205
rect -4391 1165 -4379 1199
rect -4311 1165 -4299 1199
rect -4391 1159 -4299 1165
rect -4233 1199 -4141 1205
rect -4233 1165 -4221 1199
rect -4153 1165 -4141 1199
rect -4233 1159 -4141 1165
rect -4075 1199 -3983 1205
rect -4075 1165 -4063 1199
rect -3995 1165 -3983 1199
rect -4075 1159 -3983 1165
rect -3917 1199 -3825 1205
rect -3917 1165 -3905 1199
rect -3837 1165 -3825 1199
rect -3917 1159 -3825 1165
rect -3759 1199 -3667 1205
rect -3759 1165 -3747 1199
rect -3679 1165 -3667 1199
rect -3759 1159 -3667 1165
rect -3601 1199 -3509 1205
rect -3601 1165 -3589 1199
rect -3521 1165 -3509 1199
rect -3601 1159 -3509 1165
rect -3443 1199 -3351 1205
rect -3443 1165 -3431 1199
rect -3363 1165 -3351 1199
rect -3443 1159 -3351 1165
rect -3285 1199 -3193 1205
rect -3285 1165 -3273 1199
rect -3205 1165 -3193 1199
rect -3285 1159 -3193 1165
rect -3127 1199 -3035 1205
rect -3127 1165 -3115 1199
rect -3047 1165 -3035 1199
rect -3127 1159 -3035 1165
rect -2969 1199 -2877 1205
rect -2969 1165 -2957 1199
rect -2889 1165 -2877 1199
rect -2969 1159 -2877 1165
rect -2811 1199 -2719 1205
rect -2811 1165 -2799 1199
rect -2731 1165 -2719 1199
rect -2811 1159 -2719 1165
rect -2653 1199 -2561 1205
rect -2653 1165 -2641 1199
rect -2573 1165 -2561 1199
rect -2653 1159 -2561 1165
rect -2495 1199 -2403 1205
rect -2495 1165 -2483 1199
rect -2415 1165 -2403 1199
rect -2495 1159 -2403 1165
rect -2337 1199 -2245 1205
rect -2337 1165 -2325 1199
rect -2257 1165 -2245 1199
rect -2337 1159 -2245 1165
rect -2179 1199 -2087 1205
rect -2179 1165 -2167 1199
rect -2099 1165 -2087 1199
rect -2179 1159 -2087 1165
rect -2021 1199 -1929 1205
rect -2021 1165 -2009 1199
rect -1941 1165 -1929 1199
rect -2021 1159 -1929 1165
rect -1863 1199 -1771 1205
rect -1863 1165 -1851 1199
rect -1783 1165 -1771 1199
rect -1863 1159 -1771 1165
rect -1705 1199 -1613 1205
rect -1705 1165 -1693 1199
rect -1625 1165 -1613 1199
rect -1705 1159 -1613 1165
rect -1547 1199 -1455 1205
rect -1547 1165 -1535 1199
rect -1467 1165 -1455 1199
rect -1547 1159 -1455 1165
rect -1389 1199 -1297 1205
rect -1389 1165 -1377 1199
rect -1309 1165 -1297 1199
rect -1389 1159 -1297 1165
rect -1231 1199 -1139 1205
rect -1231 1165 -1219 1199
rect -1151 1165 -1139 1199
rect -1231 1159 -1139 1165
rect -1073 1199 -981 1205
rect -1073 1165 -1061 1199
rect -993 1165 -981 1199
rect -1073 1159 -981 1165
rect -915 1199 -823 1205
rect -915 1165 -903 1199
rect -835 1165 -823 1199
rect -915 1159 -823 1165
rect -757 1199 -665 1205
rect -757 1165 -745 1199
rect -677 1165 -665 1199
rect -757 1159 -665 1165
rect -599 1199 -507 1205
rect -599 1165 -587 1199
rect -519 1165 -507 1199
rect -599 1159 -507 1165
rect -441 1199 -349 1205
rect -441 1165 -429 1199
rect -361 1165 -349 1199
rect -441 1159 -349 1165
rect -283 1199 -191 1205
rect -283 1165 -271 1199
rect -203 1165 -191 1199
rect -283 1159 -191 1165
rect -125 1199 -33 1205
rect -125 1165 -113 1199
rect -45 1165 -33 1199
rect -125 1159 -33 1165
rect 33 1199 125 1205
rect 33 1165 45 1199
rect 113 1165 125 1199
rect 33 1159 125 1165
rect 191 1199 283 1205
rect 191 1165 203 1199
rect 271 1165 283 1199
rect 191 1159 283 1165
rect 349 1199 441 1205
rect 349 1165 361 1199
rect 429 1165 441 1199
rect 349 1159 441 1165
rect 507 1199 599 1205
rect 507 1165 519 1199
rect 587 1165 599 1199
rect 507 1159 599 1165
rect 665 1199 757 1205
rect 665 1165 677 1199
rect 745 1165 757 1199
rect 665 1159 757 1165
rect 823 1199 915 1205
rect 823 1165 835 1199
rect 903 1165 915 1199
rect 823 1159 915 1165
rect 981 1199 1073 1205
rect 981 1165 993 1199
rect 1061 1165 1073 1199
rect 981 1159 1073 1165
rect 1139 1199 1231 1205
rect 1139 1165 1151 1199
rect 1219 1165 1231 1199
rect 1139 1159 1231 1165
rect 1297 1199 1389 1205
rect 1297 1165 1309 1199
rect 1377 1165 1389 1199
rect 1297 1159 1389 1165
rect 1455 1199 1547 1205
rect 1455 1165 1467 1199
rect 1535 1165 1547 1199
rect 1455 1159 1547 1165
rect 1613 1199 1705 1205
rect 1613 1165 1625 1199
rect 1693 1165 1705 1199
rect 1613 1159 1705 1165
rect 1771 1199 1863 1205
rect 1771 1165 1783 1199
rect 1851 1165 1863 1199
rect 1771 1159 1863 1165
rect 1929 1199 2021 1205
rect 1929 1165 1941 1199
rect 2009 1165 2021 1199
rect 1929 1159 2021 1165
rect 2087 1199 2179 1205
rect 2087 1165 2099 1199
rect 2167 1165 2179 1199
rect 2087 1159 2179 1165
rect 2245 1199 2337 1205
rect 2245 1165 2257 1199
rect 2325 1165 2337 1199
rect 2245 1159 2337 1165
rect 2403 1199 2495 1205
rect 2403 1165 2415 1199
rect 2483 1165 2495 1199
rect 2403 1159 2495 1165
rect 2561 1199 2653 1205
rect 2561 1165 2573 1199
rect 2641 1165 2653 1199
rect 2561 1159 2653 1165
rect 2719 1199 2811 1205
rect 2719 1165 2731 1199
rect 2799 1165 2811 1199
rect 2719 1159 2811 1165
rect 2877 1199 2969 1205
rect 2877 1165 2889 1199
rect 2957 1165 2969 1199
rect 2877 1159 2969 1165
rect 3035 1199 3127 1205
rect 3035 1165 3047 1199
rect 3115 1165 3127 1199
rect 3035 1159 3127 1165
rect 3193 1199 3285 1205
rect 3193 1165 3205 1199
rect 3273 1165 3285 1199
rect 3193 1159 3285 1165
rect 3351 1199 3443 1205
rect 3351 1165 3363 1199
rect 3431 1165 3443 1199
rect 3351 1159 3443 1165
rect 3509 1199 3601 1205
rect 3509 1165 3521 1199
rect 3589 1165 3601 1199
rect 3509 1159 3601 1165
rect 3667 1199 3759 1205
rect 3667 1165 3679 1199
rect 3747 1165 3759 1199
rect 3667 1159 3759 1165
rect 3825 1199 3917 1205
rect 3825 1165 3837 1199
rect 3905 1165 3917 1199
rect 3825 1159 3917 1165
rect 3983 1199 4075 1205
rect 3983 1165 3995 1199
rect 4063 1165 4075 1199
rect 3983 1159 4075 1165
rect 4141 1199 4233 1205
rect 4141 1165 4153 1199
rect 4221 1165 4233 1199
rect 4141 1159 4233 1165
rect 4299 1199 4391 1205
rect 4299 1165 4311 1199
rect 4379 1165 4391 1199
rect 4299 1159 4391 1165
rect 4457 1199 4549 1205
rect 4457 1165 4469 1199
rect 4537 1165 4549 1199
rect 4457 1159 4549 1165
rect 4615 1199 4707 1205
rect 4615 1165 4627 1199
rect 4695 1165 4707 1199
rect 4615 1159 4707 1165
rect 4773 1199 4865 1205
rect 4773 1165 4785 1199
rect 4853 1165 4865 1199
rect 4773 1159 4865 1165
rect -4921 1106 -4875 1118
rect -4921 130 -4915 1106
rect -4881 130 -4875 1106
rect -4921 118 -4875 130
rect -4763 1106 -4717 1118
rect -4763 130 -4757 1106
rect -4723 130 -4717 1106
rect -4763 118 -4717 130
rect -4605 1106 -4559 1118
rect -4605 130 -4599 1106
rect -4565 130 -4559 1106
rect -4605 118 -4559 130
rect -4447 1106 -4401 1118
rect -4447 130 -4441 1106
rect -4407 130 -4401 1106
rect -4447 118 -4401 130
rect -4289 1106 -4243 1118
rect -4289 130 -4283 1106
rect -4249 130 -4243 1106
rect -4289 118 -4243 130
rect -4131 1106 -4085 1118
rect -4131 130 -4125 1106
rect -4091 130 -4085 1106
rect -4131 118 -4085 130
rect -3973 1106 -3927 1118
rect -3973 130 -3967 1106
rect -3933 130 -3927 1106
rect -3973 118 -3927 130
rect -3815 1106 -3769 1118
rect -3815 130 -3809 1106
rect -3775 130 -3769 1106
rect -3815 118 -3769 130
rect -3657 1106 -3611 1118
rect -3657 130 -3651 1106
rect -3617 130 -3611 1106
rect -3657 118 -3611 130
rect -3499 1106 -3453 1118
rect -3499 130 -3493 1106
rect -3459 130 -3453 1106
rect -3499 118 -3453 130
rect -3341 1106 -3295 1118
rect -3341 130 -3335 1106
rect -3301 130 -3295 1106
rect -3341 118 -3295 130
rect -3183 1106 -3137 1118
rect -3183 130 -3177 1106
rect -3143 130 -3137 1106
rect -3183 118 -3137 130
rect -3025 1106 -2979 1118
rect -3025 130 -3019 1106
rect -2985 130 -2979 1106
rect -3025 118 -2979 130
rect -2867 1106 -2821 1118
rect -2867 130 -2861 1106
rect -2827 130 -2821 1106
rect -2867 118 -2821 130
rect -2709 1106 -2663 1118
rect -2709 130 -2703 1106
rect -2669 130 -2663 1106
rect -2709 118 -2663 130
rect -2551 1106 -2505 1118
rect -2551 130 -2545 1106
rect -2511 130 -2505 1106
rect -2551 118 -2505 130
rect -2393 1106 -2347 1118
rect -2393 130 -2387 1106
rect -2353 130 -2347 1106
rect -2393 118 -2347 130
rect -2235 1106 -2189 1118
rect -2235 130 -2229 1106
rect -2195 130 -2189 1106
rect -2235 118 -2189 130
rect -2077 1106 -2031 1118
rect -2077 130 -2071 1106
rect -2037 130 -2031 1106
rect -2077 118 -2031 130
rect -1919 1106 -1873 1118
rect -1919 130 -1913 1106
rect -1879 130 -1873 1106
rect -1919 118 -1873 130
rect -1761 1106 -1715 1118
rect -1761 130 -1755 1106
rect -1721 130 -1715 1106
rect -1761 118 -1715 130
rect -1603 1106 -1557 1118
rect -1603 130 -1597 1106
rect -1563 130 -1557 1106
rect -1603 118 -1557 130
rect -1445 1106 -1399 1118
rect -1445 130 -1439 1106
rect -1405 130 -1399 1106
rect -1445 118 -1399 130
rect -1287 1106 -1241 1118
rect -1287 130 -1281 1106
rect -1247 130 -1241 1106
rect -1287 118 -1241 130
rect -1129 1106 -1083 1118
rect -1129 130 -1123 1106
rect -1089 130 -1083 1106
rect -1129 118 -1083 130
rect -971 1106 -925 1118
rect -971 130 -965 1106
rect -931 130 -925 1106
rect -971 118 -925 130
rect -813 1106 -767 1118
rect -813 130 -807 1106
rect -773 130 -767 1106
rect -813 118 -767 130
rect -655 1106 -609 1118
rect -655 130 -649 1106
rect -615 130 -609 1106
rect -655 118 -609 130
rect -497 1106 -451 1118
rect -497 130 -491 1106
rect -457 130 -451 1106
rect -497 118 -451 130
rect -339 1106 -293 1118
rect -339 130 -333 1106
rect -299 130 -293 1106
rect -339 118 -293 130
rect -181 1106 -135 1118
rect -181 130 -175 1106
rect -141 130 -135 1106
rect -181 118 -135 130
rect -23 1106 23 1118
rect -23 130 -17 1106
rect 17 130 23 1106
rect -23 118 23 130
rect 135 1106 181 1118
rect 135 130 141 1106
rect 175 130 181 1106
rect 135 118 181 130
rect 293 1106 339 1118
rect 293 130 299 1106
rect 333 130 339 1106
rect 293 118 339 130
rect 451 1106 497 1118
rect 451 130 457 1106
rect 491 130 497 1106
rect 451 118 497 130
rect 609 1106 655 1118
rect 609 130 615 1106
rect 649 130 655 1106
rect 609 118 655 130
rect 767 1106 813 1118
rect 767 130 773 1106
rect 807 130 813 1106
rect 767 118 813 130
rect 925 1106 971 1118
rect 925 130 931 1106
rect 965 130 971 1106
rect 925 118 971 130
rect 1083 1106 1129 1118
rect 1083 130 1089 1106
rect 1123 130 1129 1106
rect 1083 118 1129 130
rect 1241 1106 1287 1118
rect 1241 130 1247 1106
rect 1281 130 1287 1106
rect 1241 118 1287 130
rect 1399 1106 1445 1118
rect 1399 130 1405 1106
rect 1439 130 1445 1106
rect 1399 118 1445 130
rect 1557 1106 1603 1118
rect 1557 130 1563 1106
rect 1597 130 1603 1106
rect 1557 118 1603 130
rect 1715 1106 1761 1118
rect 1715 130 1721 1106
rect 1755 130 1761 1106
rect 1715 118 1761 130
rect 1873 1106 1919 1118
rect 1873 130 1879 1106
rect 1913 130 1919 1106
rect 1873 118 1919 130
rect 2031 1106 2077 1118
rect 2031 130 2037 1106
rect 2071 130 2077 1106
rect 2031 118 2077 130
rect 2189 1106 2235 1118
rect 2189 130 2195 1106
rect 2229 130 2235 1106
rect 2189 118 2235 130
rect 2347 1106 2393 1118
rect 2347 130 2353 1106
rect 2387 130 2393 1106
rect 2347 118 2393 130
rect 2505 1106 2551 1118
rect 2505 130 2511 1106
rect 2545 130 2551 1106
rect 2505 118 2551 130
rect 2663 1106 2709 1118
rect 2663 130 2669 1106
rect 2703 130 2709 1106
rect 2663 118 2709 130
rect 2821 1106 2867 1118
rect 2821 130 2827 1106
rect 2861 130 2867 1106
rect 2821 118 2867 130
rect 2979 1106 3025 1118
rect 2979 130 2985 1106
rect 3019 130 3025 1106
rect 2979 118 3025 130
rect 3137 1106 3183 1118
rect 3137 130 3143 1106
rect 3177 130 3183 1106
rect 3137 118 3183 130
rect 3295 1106 3341 1118
rect 3295 130 3301 1106
rect 3335 130 3341 1106
rect 3295 118 3341 130
rect 3453 1106 3499 1118
rect 3453 130 3459 1106
rect 3493 130 3499 1106
rect 3453 118 3499 130
rect 3611 1106 3657 1118
rect 3611 130 3617 1106
rect 3651 130 3657 1106
rect 3611 118 3657 130
rect 3769 1106 3815 1118
rect 3769 130 3775 1106
rect 3809 130 3815 1106
rect 3769 118 3815 130
rect 3927 1106 3973 1118
rect 3927 130 3933 1106
rect 3967 130 3973 1106
rect 3927 118 3973 130
rect 4085 1106 4131 1118
rect 4085 130 4091 1106
rect 4125 130 4131 1106
rect 4085 118 4131 130
rect 4243 1106 4289 1118
rect 4243 130 4249 1106
rect 4283 130 4289 1106
rect 4243 118 4289 130
rect 4401 1106 4447 1118
rect 4401 130 4407 1106
rect 4441 130 4447 1106
rect 4401 118 4447 130
rect 4559 1106 4605 1118
rect 4559 130 4565 1106
rect 4599 130 4605 1106
rect 4559 118 4605 130
rect 4717 1106 4763 1118
rect 4717 130 4723 1106
rect 4757 130 4763 1106
rect 4717 118 4763 130
rect 4875 1106 4921 1118
rect 4875 130 4881 1106
rect 4915 130 4921 1106
rect 4875 118 4921 130
rect -4865 71 -4773 77
rect -4865 37 -4853 71
rect -4785 37 -4773 71
rect -4865 31 -4773 37
rect -4707 71 -4615 77
rect -4707 37 -4695 71
rect -4627 37 -4615 71
rect -4707 31 -4615 37
rect -4549 71 -4457 77
rect -4549 37 -4537 71
rect -4469 37 -4457 71
rect -4549 31 -4457 37
rect -4391 71 -4299 77
rect -4391 37 -4379 71
rect -4311 37 -4299 71
rect -4391 31 -4299 37
rect -4233 71 -4141 77
rect -4233 37 -4221 71
rect -4153 37 -4141 71
rect -4233 31 -4141 37
rect -4075 71 -3983 77
rect -4075 37 -4063 71
rect -3995 37 -3983 71
rect -4075 31 -3983 37
rect -3917 71 -3825 77
rect -3917 37 -3905 71
rect -3837 37 -3825 71
rect -3917 31 -3825 37
rect -3759 71 -3667 77
rect -3759 37 -3747 71
rect -3679 37 -3667 71
rect -3759 31 -3667 37
rect -3601 71 -3509 77
rect -3601 37 -3589 71
rect -3521 37 -3509 71
rect -3601 31 -3509 37
rect -3443 71 -3351 77
rect -3443 37 -3431 71
rect -3363 37 -3351 71
rect -3443 31 -3351 37
rect -3285 71 -3193 77
rect -3285 37 -3273 71
rect -3205 37 -3193 71
rect -3285 31 -3193 37
rect -3127 71 -3035 77
rect -3127 37 -3115 71
rect -3047 37 -3035 71
rect -3127 31 -3035 37
rect -2969 71 -2877 77
rect -2969 37 -2957 71
rect -2889 37 -2877 71
rect -2969 31 -2877 37
rect -2811 71 -2719 77
rect -2811 37 -2799 71
rect -2731 37 -2719 71
rect -2811 31 -2719 37
rect -2653 71 -2561 77
rect -2653 37 -2641 71
rect -2573 37 -2561 71
rect -2653 31 -2561 37
rect -2495 71 -2403 77
rect -2495 37 -2483 71
rect -2415 37 -2403 71
rect -2495 31 -2403 37
rect -2337 71 -2245 77
rect -2337 37 -2325 71
rect -2257 37 -2245 71
rect -2337 31 -2245 37
rect -2179 71 -2087 77
rect -2179 37 -2167 71
rect -2099 37 -2087 71
rect -2179 31 -2087 37
rect -2021 71 -1929 77
rect -2021 37 -2009 71
rect -1941 37 -1929 71
rect -2021 31 -1929 37
rect -1863 71 -1771 77
rect -1863 37 -1851 71
rect -1783 37 -1771 71
rect -1863 31 -1771 37
rect -1705 71 -1613 77
rect -1705 37 -1693 71
rect -1625 37 -1613 71
rect -1705 31 -1613 37
rect -1547 71 -1455 77
rect -1547 37 -1535 71
rect -1467 37 -1455 71
rect -1547 31 -1455 37
rect -1389 71 -1297 77
rect -1389 37 -1377 71
rect -1309 37 -1297 71
rect -1389 31 -1297 37
rect -1231 71 -1139 77
rect -1231 37 -1219 71
rect -1151 37 -1139 71
rect -1231 31 -1139 37
rect -1073 71 -981 77
rect -1073 37 -1061 71
rect -993 37 -981 71
rect -1073 31 -981 37
rect -915 71 -823 77
rect -915 37 -903 71
rect -835 37 -823 71
rect -915 31 -823 37
rect -757 71 -665 77
rect -757 37 -745 71
rect -677 37 -665 71
rect -757 31 -665 37
rect -599 71 -507 77
rect -599 37 -587 71
rect -519 37 -507 71
rect -599 31 -507 37
rect -441 71 -349 77
rect -441 37 -429 71
rect -361 37 -349 71
rect -441 31 -349 37
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect 349 71 441 77
rect 349 37 361 71
rect 429 37 441 71
rect 349 31 441 37
rect 507 71 599 77
rect 507 37 519 71
rect 587 37 599 71
rect 507 31 599 37
rect 665 71 757 77
rect 665 37 677 71
rect 745 37 757 71
rect 665 31 757 37
rect 823 71 915 77
rect 823 37 835 71
rect 903 37 915 71
rect 823 31 915 37
rect 981 71 1073 77
rect 981 37 993 71
rect 1061 37 1073 71
rect 981 31 1073 37
rect 1139 71 1231 77
rect 1139 37 1151 71
rect 1219 37 1231 71
rect 1139 31 1231 37
rect 1297 71 1389 77
rect 1297 37 1309 71
rect 1377 37 1389 71
rect 1297 31 1389 37
rect 1455 71 1547 77
rect 1455 37 1467 71
rect 1535 37 1547 71
rect 1455 31 1547 37
rect 1613 71 1705 77
rect 1613 37 1625 71
rect 1693 37 1705 71
rect 1613 31 1705 37
rect 1771 71 1863 77
rect 1771 37 1783 71
rect 1851 37 1863 71
rect 1771 31 1863 37
rect 1929 71 2021 77
rect 1929 37 1941 71
rect 2009 37 2021 71
rect 1929 31 2021 37
rect 2087 71 2179 77
rect 2087 37 2099 71
rect 2167 37 2179 71
rect 2087 31 2179 37
rect 2245 71 2337 77
rect 2245 37 2257 71
rect 2325 37 2337 71
rect 2245 31 2337 37
rect 2403 71 2495 77
rect 2403 37 2415 71
rect 2483 37 2495 71
rect 2403 31 2495 37
rect 2561 71 2653 77
rect 2561 37 2573 71
rect 2641 37 2653 71
rect 2561 31 2653 37
rect 2719 71 2811 77
rect 2719 37 2731 71
rect 2799 37 2811 71
rect 2719 31 2811 37
rect 2877 71 2969 77
rect 2877 37 2889 71
rect 2957 37 2969 71
rect 2877 31 2969 37
rect 3035 71 3127 77
rect 3035 37 3047 71
rect 3115 37 3127 71
rect 3035 31 3127 37
rect 3193 71 3285 77
rect 3193 37 3205 71
rect 3273 37 3285 71
rect 3193 31 3285 37
rect 3351 71 3443 77
rect 3351 37 3363 71
rect 3431 37 3443 71
rect 3351 31 3443 37
rect 3509 71 3601 77
rect 3509 37 3521 71
rect 3589 37 3601 71
rect 3509 31 3601 37
rect 3667 71 3759 77
rect 3667 37 3679 71
rect 3747 37 3759 71
rect 3667 31 3759 37
rect 3825 71 3917 77
rect 3825 37 3837 71
rect 3905 37 3917 71
rect 3825 31 3917 37
rect 3983 71 4075 77
rect 3983 37 3995 71
rect 4063 37 4075 71
rect 3983 31 4075 37
rect 4141 71 4233 77
rect 4141 37 4153 71
rect 4221 37 4233 71
rect 4141 31 4233 37
rect 4299 71 4391 77
rect 4299 37 4311 71
rect 4379 37 4391 71
rect 4299 31 4391 37
rect 4457 71 4549 77
rect 4457 37 4469 71
rect 4537 37 4549 71
rect 4457 31 4549 37
rect 4615 71 4707 77
rect 4615 37 4627 71
rect 4695 37 4707 71
rect 4615 31 4707 37
rect 4773 71 4865 77
rect 4773 37 4785 71
rect 4853 37 4865 71
rect 4773 31 4865 37
rect -4865 -37 -4773 -31
rect -4865 -71 -4853 -37
rect -4785 -71 -4773 -37
rect -4865 -77 -4773 -71
rect -4707 -37 -4615 -31
rect -4707 -71 -4695 -37
rect -4627 -71 -4615 -37
rect -4707 -77 -4615 -71
rect -4549 -37 -4457 -31
rect -4549 -71 -4537 -37
rect -4469 -71 -4457 -37
rect -4549 -77 -4457 -71
rect -4391 -37 -4299 -31
rect -4391 -71 -4379 -37
rect -4311 -71 -4299 -37
rect -4391 -77 -4299 -71
rect -4233 -37 -4141 -31
rect -4233 -71 -4221 -37
rect -4153 -71 -4141 -37
rect -4233 -77 -4141 -71
rect -4075 -37 -3983 -31
rect -4075 -71 -4063 -37
rect -3995 -71 -3983 -37
rect -4075 -77 -3983 -71
rect -3917 -37 -3825 -31
rect -3917 -71 -3905 -37
rect -3837 -71 -3825 -37
rect -3917 -77 -3825 -71
rect -3759 -37 -3667 -31
rect -3759 -71 -3747 -37
rect -3679 -71 -3667 -37
rect -3759 -77 -3667 -71
rect -3601 -37 -3509 -31
rect -3601 -71 -3589 -37
rect -3521 -71 -3509 -37
rect -3601 -77 -3509 -71
rect -3443 -37 -3351 -31
rect -3443 -71 -3431 -37
rect -3363 -71 -3351 -37
rect -3443 -77 -3351 -71
rect -3285 -37 -3193 -31
rect -3285 -71 -3273 -37
rect -3205 -71 -3193 -37
rect -3285 -77 -3193 -71
rect -3127 -37 -3035 -31
rect -3127 -71 -3115 -37
rect -3047 -71 -3035 -37
rect -3127 -77 -3035 -71
rect -2969 -37 -2877 -31
rect -2969 -71 -2957 -37
rect -2889 -71 -2877 -37
rect -2969 -77 -2877 -71
rect -2811 -37 -2719 -31
rect -2811 -71 -2799 -37
rect -2731 -71 -2719 -37
rect -2811 -77 -2719 -71
rect -2653 -37 -2561 -31
rect -2653 -71 -2641 -37
rect -2573 -71 -2561 -37
rect -2653 -77 -2561 -71
rect -2495 -37 -2403 -31
rect -2495 -71 -2483 -37
rect -2415 -71 -2403 -37
rect -2495 -77 -2403 -71
rect -2337 -37 -2245 -31
rect -2337 -71 -2325 -37
rect -2257 -71 -2245 -37
rect -2337 -77 -2245 -71
rect -2179 -37 -2087 -31
rect -2179 -71 -2167 -37
rect -2099 -71 -2087 -37
rect -2179 -77 -2087 -71
rect -2021 -37 -1929 -31
rect -2021 -71 -2009 -37
rect -1941 -71 -1929 -37
rect -2021 -77 -1929 -71
rect -1863 -37 -1771 -31
rect -1863 -71 -1851 -37
rect -1783 -71 -1771 -37
rect -1863 -77 -1771 -71
rect -1705 -37 -1613 -31
rect -1705 -71 -1693 -37
rect -1625 -71 -1613 -37
rect -1705 -77 -1613 -71
rect -1547 -37 -1455 -31
rect -1547 -71 -1535 -37
rect -1467 -71 -1455 -37
rect -1547 -77 -1455 -71
rect -1389 -37 -1297 -31
rect -1389 -71 -1377 -37
rect -1309 -71 -1297 -37
rect -1389 -77 -1297 -71
rect -1231 -37 -1139 -31
rect -1231 -71 -1219 -37
rect -1151 -71 -1139 -37
rect -1231 -77 -1139 -71
rect -1073 -37 -981 -31
rect -1073 -71 -1061 -37
rect -993 -71 -981 -37
rect -1073 -77 -981 -71
rect -915 -37 -823 -31
rect -915 -71 -903 -37
rect -835 -71 -823 -37
rect -915 -77 -823 -71
rect -757 -37 -665 -31
rect -757 -71 -745 -37
rect -677 -71 -665 -37
rect -757 -77 -665 -71
rect -599 -37 -507 -31
rect -599 -71 -587 -37
rect -519 -71 -507 -37
rect -599 -77 -507 -71
rect -441 -37 -349 -31
rect -441 -71 -429 -37
rect -361 -71 -349 -37
rect -441 -77 -349 -71
rect -283 -37 -191 -31
rect -283 -71 -271 -37
rect -203 -71 -191 -37
rect -283 -77 -191 -71
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect 191 -37 283 -31
rect 191 -71 203 -37
rect 271 -71 283 -37
rect 191 -77 283 -71
rect 349 -37 441 -31
rect 349 -71 361 -37
rect 429 -71 441 -37
rect 349 -77 441 -71
rect 507 -37 599 -31
rect 507 -71 519 -37
rect 587 -71 599 -37
rect 507 -77 599 -71
rect 665 -37 757 -31
rect 665 -71 677 -37
rect 745 -71 757 -37
rect 665 -77 757 -71
rect 823 -37 915 -31
rect 823 -71 835 -37
rect 903 -71 915 -37
rect 823 -77 915 -71
rect 981 -37 1073 -31
rect 981 -71 993 -37
rect 1061 -71 1073 -37
rect 981 -77 1073 -71
rect 1139 -37 1231 -31
rect 1139 -71 1151 -37
rect 1219 -71 1231 -37
rect 1139 -77 1231 -71
rect 1297 -37 1389 -31
rect 1297 -71 1309 -37
rect 1377 -71 1389 -37
rect 1297 -77 1389 -71
rect 1455 -37 1547 -31
rect 1455 -71 1467 -37
rect 1535 -71 1547 -37
rect 1455 -77 1547 -71
rect 1613 -37 1705 -31
rect 1613 -71 1625 -37
rect 1693 -71 1705 -37
rect 1613 -77 1705 -71
rect 1771 -37 1863 -31
rect 1771 -71 1783 -37
rect 1851 -71 1863 -37
rect 1771 -77 1863 -71
rect 1929 -37 2021 -31
rect 1929 -71 1941 -37
rect 2009 -71 2021 -37
rect 1929 -77 2021 -71
rect 2087 -37 2179 -31
rect 2087 -71 2099 -37
rect 2167 -71 2179 -37
rect 2087 -77 2179 -71
rect 2245 -37 2337 -31
rect 2245 -71 2257 -37
rect 2325 -71 2337 -37
rect 2245 -77 2337 -71
rect 2403 -37 2495 -31
rect 2403 -71 2415 -37
rect 2483 -71 2495 -37
rect 2403 -77 2495 -71
rect 2561 -37 2653 -31
rect 2561 -71 2573 -37
rect 2641 -71 2653 -37
rect 2561 -77 2653 -71
rect 2719 -37 2811 -31
rect 2719 -71 2731 -37
rect 2799 -71 2811 -37
rect 2719 -77 2811 -71
rect 2877 -37 2969 -31
rect 2877 -71 2889 -37
rect 2957 -71 2969 -37
rect 2877 -77 2969 -71
rect 3035 -37 3127 -31
rect 3035 -71 3047 -37
rect 3115 -71 3127 -37
rect 3035 -77 3127 -71
rect 3193 -37 3285 -31
rect 3193 -71 3205 -37
rect 3273 -71 3285 -37
rect 3193 -77 3285 -71
rect 3351 -37 3443 -31
rect 3351 -71 3363 -37
rect 3431 -71 3443 -37
rect 3351 -77 3443 -71
rect 3509 -37 3601 -31
rect 3509 -71 3521 -37
rect 3589 -71 3601 -37
rect 3509 -77 3601 -71
rect 3667 -37 3759 -31
rect 3667 -71 3679 -37
rect 3747 -71 3759 -37
rect 3667 -77 3759 -71
rect 3825 -37 3917 -31
rect 3825 -71 3837 -37
rect 3905 -71 3917 -37
rect 3825 -77 3917 -71
rect 3983 -37 4075 -31
rect 3983 -71 3995 -37
rect 4063 -71 4075 -37
rect 3983 -77 4075 -71
rect 4141 -37 4233 -31
rect 4141 -71 4153 -37
rect 4221 -71 4233 -37
rect 4141 -77 4233 -71
rect 4299 -37 4391 -31
rect 4299 -71 4311 -37
rect 4379 -71 4391 -37
rect 4299 -77 4391 -71
rect 4457 -37 4549 -31
rect 4457 -71 4469 -37
rect 4537 -71 4549 -37
rect 4457 -77 4549 -71
rect 4615 -37 4707 -31
rect 4615 -71 4627 -37
rect 4695 -71 4707 -37
rect 4615 -77 4707 -71
rect 4773 -37 4865 -31
rect 4773 -71 4785 -37
rect 4853 -71 4865 -37
rect 4773 -77 4865 -71
rect -4921 -130 -4875 -118
rect -4921 -1106 -4915 -130
rect -4881 -1106 -4875 -130
rect -4921 -1118 -4875 -1106
rect -4763 -130 -4717 -118
rect -4763 -1106 -4757 -130
rect -4723 -1106 -4717 -130
rect -4763 -1118 -4717 -1106
rect -4605 -130 -4559 -118
rect -4605 -1106 -4599 -130
rect -4565 -1106 -4559 -130
rect -4605 -1118 -4559 -1106
rect -4447 -130 -4401 -118
rect -4447 -1106 -4441 -130
rect -4407 -1106 -4401 -130
rect -4447 -1118 -4401 -1106
rect -4289 -130 -4243 -118
rect -4289 -1106 -4283 -130
rect -4249 -1106 -4243 -130
rect -4289 -1118 -4243 -1106
rect -4131 -130 -4085 -118
rect -4131 -1106 -4125 -130
rect -4091 -1106 -4085 -130
rect -4131 -1118 -4085 -1106
rect -3973 -130 -3927 -118
rect -3973 -1106 -3967 -130
rect -3933 -1106 -3927 -130
rect -3973 -1118 -3927 -1106
rect -3815 -130 -3769 -118
rect -3815 -1106 -3809 -130
rect -3775 -1106 -3769 -130
rect -3815 -1118 -3769 -1106
rect -3657 -130 -3611 -118
rect -3657 -1106 -3651 -130
rect -3617 -1106 -3611 -130
rect -3657 -1118 -3611 -1106
rect -3499 -130 -3453 -118
rect -3499 -1106 -3493 -130
rect -3459 -1106 -3453 -130
rect -3499 -1118 -3453 -1106
rect -3341 -130 -3295 -118
rect -3341 -1106 -3335 -130
rect -3301 -1106 -3295 -130
rect -3341 -1118 -3295 -1106
rect -3183 -130 -3137 -118
rect -3183 -1106 -3177 -130
rect -3143 -1106 -3137 -130
rect -3183 -1118 -3137 -1106
rect -3025 -130 -2979 -118
rect -3025 -1106 -3019 -130
rect -2985 -1106 -2979 -130
rect -3025 -1118 -2979 -1106
rect -2867 -130 -2821 -118
rect -2867 -1106 -2861 -130
rect -2827 -1106 -2821 -130
rect -2867 -1118 -2821 -1106
rect -2709 -130 -2663 -118
rect -2709 -1106 -2703 -130
rect -2669 -1106 -2663 -130
rect -2709 -1118 -2663 -1106
rect -2551 -130 -2505 -118
rect -2551 -1106 -2545 -130
rect -2511 -1106 -2505 -130
rect -2551 -1118 -2505 -1106
rect -2393 -130 -2347 -118
rect -2393 -1106 -2387 -130
rect -2353 -1106 -2347 -130
rect -2393 -1118 -2347 -1106
rect -2235 -130 -2189 -118
rect -2235 -1106 -2229 -130
rect -2195 -1106 -2189 -130
rect -2235 -1118 -2189 -1106
rect -2077 -130 -2031 -118
rect -2077 -1106 -2071 -130
rect -2037 -1106 -2031 -130
rect -2077 -1118 -2031 -1106
rect -1919 -130 -1873 -118
rect -1919 -1106 -1913 -130
rect -1879 -1106 -1873 -130
rect -1919 -1118 -1873 -1106
rect -1761 -130 -1715 -118
rect -1761 -1106 -1755 -130
rect -1721 -1106 -1715 -130
rect -1761 -1118 -1715 -1106
rect -1603 -130 -1557 -118
rect -1603 -1106 -1597 -130
rect -1563 -1106 -1557 -130
rect -1603 -1118 -1557 -1106
rect -1445 -130 -1399 -118
rect -1445 -1106 -1439 -130
rect -1405 -1106 -1399 -130
rect -1445 -1118 -1399 -1106
rect -1287 -130 -1241 -118
rect -1287 -1106 -1281 -130
rect -1247 -1106 -1241 -130
rect -1287 -1118 -1241 -1106
rect -1129 -130 -1083 -118
rect -1129 -1106 -1123 -130
rect -1089 -1106 -1083 -130
rect -1129 -1118 -1083 -1106
rect -971 -130 -925 -118
rect -971 -1106 -965 -130
rect -931 -1106 -925 -130
rect -971 -1118 -925 -1106
rect -813 -130 -767 -118
rect -813 -1106 -807 -130
rect -773 -1106 -767 -130
rect -813 -1118 -767 -1106
rect -655 -130 -609 -118
rect -655 -1106 -649 -130
rect -615 -1106 -609 -130
rect -655 -1118 -609 -1106
rect -497 -130 -451 -118
rect -497 -1106 -491 -130
rect -457 -1106 -451 -130
rect -497 -1118 -451 -1106
rect -339 -130 -293 -118
rect -339 -1106 -333 -130
rect -299 -1106 -293 -130
rect -339 -1118 -293 -1106
rect -181 -130 -135 -118
rect -181 -1106 -175 -130
rect -141 -1106 -135 -130
rect -181 -1118 -135 -1106
rect -23 -130 23 -118
rect -23 -1106 -17 -130
rect 17 -1106 23 -130
rect -23 -1118 23 -1106
rect 135 -130 181 -118
rect 135 -1106 141 -130
rect 175 -1106 181 -130
rect 135 -1118 181 -1106
rect 293 -130 339 -118
rect 293 -1106 299 -130
rect 333 -1106 339 -130
rect 293 -1118 339 -1106
rect 451 -130 497 -118
rect 451 -1106 457 -130
rect 491 -1106 497 -130
rect 451 -1118 497 -1106
rect 609 -130 655 -118
rect 609 -1106 615 -130
rect 649 -1106 655 -130
rect 609 -1118 655 -1106
rect 767 -130 813 -118
rect 767 -1106 773 -130
rect 807 -1106 813 -130
rect 767 -1118 813 -1106
rect 925 -130 971 -118
rect 925 -1106 931 -130
rect 965 -1106 971 -130
rect 925 -1118 971 -1106
rect 1083 -130 1129 -118
rect 1083 -1106 1089 -130
rect 1123 -1106 1129 -130
rect 1083 -1118 1129 -1106
rect 1241 -130 1287 -118
rect 1241 -1106 1247 -130
rect 1281 -1106 1287 -130
rect 1241 -1118 1287 -1106
rect 1399 -130 1445 -118
rect 1399 -1106 1405 -130
rect 1439 -1106 1445 -130
rect 1399 -1118 1445 -1106
rect 1557 -130 1603 -118
rect 1557 -1106 1563 -130
rect 1597 -1106 1603 -130
rect 1557 -1118 1603 -1106
rect 1715 -130 1761 -118
rect 1715 -1106 1721 -130
rect 1755 -1106 1761 -130
rect 1715 -1118 1761 -1106
rect 1873 -130 1919 -118
rect 1873 -1106 1879 -130
rect 1913 -1106 1919 -130
rect 1873 -1118 1919 -1106
rect 2031 -130 2077 -118
rect 2031 -1106 2037 -130
rect 2071 -1106 2077 -130
rect 2031 -1118 2077 -1106
rect 2189 -130 2235 -118
rect 2189 -1106 2195 -130
rect 2229 -1106 2235 -130
rect 2189 -1118 2235 -1106
rect 2347 -130 2393 -118
rect 2347 -1106 2353 -130
rect 2387 -1106 2393 -130
rect 2347 -1118 2393 -1106
rect 2505 -130 2551 -118
rect 2505 -1106 2511 -130
rect 2545 -1106 2551 -130
rect 2505 -1118 2551 -1106
rect 2663 -130 2709 -118
rect 2663 -1106 2669 -130
rect 2703 -1106 2709 -130
rect 2663 -1118 2709 -1106
rect 2821 -130 2867 -118
rect 2821 -1106 2827 -130
rect 2861 -1106 2867 -130
rect 2821 -1118 2867 -1106
rect 2979 -130 3025 -118
rect 2979 -1106 2985 -130
rect 3019 -1106 3025 -130
rect 2979 -1118 3025 -1106
rect 3137 -130 3183 -118
rect 3137 -1106 3143 -130
rect 3177 -1106 3183 -130
rect 3137 -1118 3183 -1106
rect 3295 -130 3341 -118
rect 3295 -1106 3301 -130
rect 3335 -1106 3341 -130
rect 3295 -1118 3341 -1106
rect 3453 -130 3499 -118
rect 3453 -1106 3459 -130
rect 3493 -1106 3499 -130
rect 3453 -1118 3499 -1106
rect 3611 -130 3657 -118
rect 3611 -1106 3617 -130
rect 3651 -1106 3657 -130
rect 3611 -1118 3657 -1106
rect 3769 -130 3815 -118
rect 3769 -1106 3775 -130
rect 3809 -1106 3815 -130
rect 3769 -1118 3815 -1106
rect 3927 -130 3973 -118
rect 3927 -1106 3933 -130
rect 3967 -1106 3973 -130
rect 3927 -1118 3973 -1106
rect 4085 -130 4131 -118
rect 4085 -1106 4091 -130
rect 4125 -1106 4131 -130
rect 4085 -1118 4131 -1106
rect 4243 -130 4289 -118
rect 4243 -1106 4249 -130
rect 4283 -1106 4289 -130
rect 4243 -1118 4289 -1106
rect 4401 -130 4447 -118
rect 4401 -1106 4407 -130
rect 4441 -1106 4447 -130
rect 4401 -1118 4447 -1106
rect 4559 -130 4605 -118
rect 4559 -1106 4565 -130
rect 4599 -1106 4605 -130
rect 4559 -1118 4605 -1106
rect 4717 -130 4763 -118
rect 4717 -1106 4723 -130
rect 4757 -1106 4763 -130
rect 4717 -1118 4763 -1106
rect 4875 -130 4921 -118
rect 4875 -1106 4881 -130
rect 4915 -1106 4921 -130
rect 4875 -1118 4921 -1106
rect -4865 -1165 -4773 -1159
rect -4865 -1199 -4853 -1165
rect -4785 -1199 -4773 -1165
rect -4865 -1205 -4773 -1199
rect -4707 -1165 -4615 -1159
rect -4707 -1199 -4695 -1165
rect -4627 -1199 -4615 -1165
rect -4707 -1205 -4615 -1199
rect -4549 -1165 -4457 -1159
rect -4549 -1199 -4537 -1165
rect -4469 -1199 -4457 -1165
rect -4549 -1205 -4457 -1199
rect -4391 -1165 -4299 -1159
rect -4391 -1199 -4379 -1165
rect -4311 -1199 -4299 -1165
rect -4391 -1205 -4299 -1199
rect -4233 -1165 -4141 -1159
rect -4233 -1199 -4221 -1165
rect -4153 -1199 -4141 -1165
rect -4233 -1205 -4141 -1199
rect -4075 -1165 -3983 -1159
rect -4075 -1199 -4063 -1165
rect -3995 -1199 -3983 -1165
rect -4075 -1205 -3983 -1199
rect -3917 -1165 -3825 -1159
rect -3917 -1199 -3905 -1165
rect -3837 -1199 -3825 -1165
rect -3917 -1205 -3825 -1199
rect -3759 -1165 -3667 -1159
rect -3759 -1199 -3747 -1165
rect -3679 -1199 -3667 -1165
rect -3759 -1205 -3667 -1199
rect -3601 -1165 -3509 -1159
rect -3601 -1199 -3589 -1165
rect -3521 -1199 -3509 -1165
rect -3601 -1205 -3509 -1199
rect -3443 -1165 -3351 -1159
rect -3443 -1199 -3431 -1165
rect -3363 -1199 -3351 -1165
rect -3443 -1205 -3351 -1199
rect -3285 -1165 -3193 -1159
rect -3285 -1199 -3273 -1165
rect -3205 -1199 -3193 -1165
rect -3285 -1205 -3193 -1199
rect -3127 -1165 -3035 -1159
rect -3127 -1199 -3115 -1165
rect -3047 -1199 -3035 -1165
rect -3127 -1205 -3035 -1199
rect -2969 -1165 -2877 -1159
rect -2969 -1199 -2957 -1165
rect -2889 -1199 -2877 -1165
rect -2969 -1205 -2877 -1199
rect -2811 -1165 -2719 -1159
rect -2811 -1199 -2799 -1165
rect -2731 -1199 -2719 -1165
rect -2811 -1205 -2719 -1199
rect -2653 -1165 -2561 -1159
rect -2653 -1199 -2641 -1165
rect -2573 -1199 -2561 -1165
rect -2653 -1205 -2561 -1199
rect -2495 -1165 -2403 -1159
rect -2495 -1199 -2483 -1165
rect -2415 -1199 -2403 -1165
rect -2495 -1205 -2403 -1199
rect -2337 -1165 -2245 -1159
rect -2337 -1199 -2325 -1165
rect -2257 -1199 -2245 -1165
rect -2337 -1205 -2245 -1199
rect -2179 -1165 -2087 -1159
rect -2179 -1199 -2167 -1165
rect -2099 -1199 -2087 -1165
rect -2179 -1205 -2087 -1199
rect -2021 -1165 -1929 -1159
rect -2021 -1199 -2009 -1165
rect -1941 -1199 -1929 -1165
rect -2021 -1205 -1929 -1199
rect -1863 -1165 -1771 -1159
rect -1863 -1199 -1851 -1165
rect -1783 -1199 -1771 -1165
rect -1863 -1205 -1771 -1199
rect -1705 -1165 -1613 -1159
rect -1705 -1199 -1693 -1165
rect -1625 -1199 -1613 -1165
rect -1705 -1205 -1613 -1199
rect -1547 -1165 -1455 -1159
rect -1547 -1199 -1535 -1165
rect -1467 -1199 -1455 -1165
rect -1547 -1205 -1455 -1199
rect -1389 -1165 -1297 -1159
rect -1389 -1199 -1377 -1165
rect -1309 -1199 -1297 -1165
rect -1389 -1205 -1297 -1199
rect -1231 -1165 -1139 -1159
rect -1231 -1199 -1219 -1165
rect -1151 -1199 -1139 -1165
rect -1231 -1205 -1139 -1199
rect -1073 -1165 -981 -1159
rect -1073 -1199 -1061 -1165
rect -993 -1199 -981 -1165
rect -1073 -1205 -981 -1199
rect -915 -1165 -823 -1159
rect -915 -1199 -903 -1165
rect -835 -1199 -823 -1165
rect -915 -1205 -823 -1199
rect -757 -1165 -665 -1159
rect -757 -1199 -745 -1165
rect -677 -1199 -665 -1165
rect -757 -1205 -665 -1199
rect -599 -1165 -507 -1159
rect -599 -1199 -587 -1165
rect -519 -1199 -507 -1165
rect -599 -1205 -507 -1199
rect -441 -1165 -349 -1159
rect -441 -1199 -429 -1165
rect -361 -1199 -349 -1165
rect -441 -1205 -349 -1199
rect -283 -1165 -191 -1159
rect -283 -1199 -271 -1165
rect -203 -1199 -191 -1165
rect -283 -1205 -191 -1199
rect -125 -1165 -33 -1159
rect -125 -1199 -113 -1165
rect -45 -1199 -33 -1165
rect -125 -1205 -33 -1199
rect 33 -1165 125 -1159
rect 33 -1199 45 -1165
rect 113 -1199 125 -1165
rect 33 -1205 125 -1199
rect 191 -1165 283 -1159
rect 191 -1199 203 -1165
rect 271 -1199 283 -1165
rect 191 -1205 283 -1199
rect 349 -1165 441 -1159
rect 349 -1199 361 -1165
rect 429 -1199 441 -1165
rect 349 -1205 441 -1199
rect 507 -1165 599 -1159
rect 507 -1199 519 -1165
rect 587 -1199 599 -1165
rect 507 -1205 599 -1199
rect 665 -1165 757 -1159
rect 665 -1199 677 -1165
rect 745 -1199 757 -1165
rect 665 -1205 757 -1199
rect 823 -1165 915 -1159
rect 823 -1199 835 -1165
rect 903 -1199 915 -1165
rect 823 -1205 915 -1199
rect 981 -1165 1073 -1159
rect 981 -1199 993 -1165
rect 1061 -1199 1073 -1165
rect 981 -1205 1073 -1199
rect 1139 -1165 1231 -1159
rect 1139 -1199 1151 -1165
rect 1219 -1199 1231 -1165
rect 1139 -1205 1231 -1199
rect 1297 -1165 1389 -1159
rect 1297 -1199 1309 -1165
rect 1377 -1199 1389 -1165
rect 1297 -1205 1389 -1199
rect 1455 -1165 1547 -1159
rect 1455 -1199 1467 -1165
rect 1535 -1199 1547 -1165
rect 1455 -1205 1547 -1199
rect 1613 -1165 1705 -1159
rect 1613 -1199 1625 -1165
rect 1693 -1199 1705 -1165
rect 1613 -1205 1705 -1199
rect 1771 -1165 1863 -1159
rect 1771 -1199 1783 -1165
rect 1851 -1199 1863 -1165
rect 1771 -1205 1863 -1199
rect 1929 -1165 2021 -1159
rect 1929 -1199 1941 -1165
rect 2009 -1199 2021 -1165
rect 1929 -1205 2021 -1199
rect 2087 -1165 2179 -1159
rect 2087 -1199 2099 -1165
rect 2167 -1199 2179 -1165
rect 2087 -1205 2179 -1199
rect 2245 -1165 2337 -1159
rect 2245 -1199 2257 -1165
rect 2325 -1199 2337 -1165
rect 2245 -1205 2337 -1199
rect 2403 -1165 2495 -1159
rect 2403 -1199 2415 -1165
rect 2483 -1199 2495 -1165
rect 2403 -1205 2495 -1199
rect 2561 -1165 2653 -1159
rect 2561 -1199 2573 -1165
rect 2641 -1199 2653 -1165
rect 2561 -1205 2653 -1199
rect 2719 -1165 2811 -1159
rect 2719 -1199 2731 -1165
rect 2799 -1199 2811 -1165
rect 2719 -1205 2811 -1199
rect 2877 -1165 2969 -1159
rect 2877 -1199 2889 -1165
rect 2957 -1199 2969 -1165
rect 2877 -1205 2969 -1199
rect 3035 -1165 3127 -1159
rect 3035 -1199 3047 -1165
rect 3115 -1199 3127 -1165
rect 3035 -1205 3127 -1199
rect 3193 -1165 3285 -1159
rect 3193 -1199 3205 -1165
rect 3273 -1199 3285 -1165
rect 3193 -1205 3285 -1199
rect 3351 -1165 3443 -1159
rect 3351 -1199 3363 -1165
rect 3431 -1199 3443 -1165
rect 3351 -1205 3443 -1199
rect 3509 -1165 3601 -1159
rect 3509 -1199 3521 -1165
rect 3589 -1199 3601 -1165
rect 3509 -1205 3601 -1199
rect 3667 -1165 3759 -1159
rect 3667 -1199 3679 -1165
rect 3747 -1199 3759 -1165
rect 3667 -1205 3759 -1199
rect 3825 -1165 3917 -1159
rect 3825 -1199 3837 -1165
rect 3905 -1199 3917 -1165
rect 3825 -1205 3917 -1199
rect 3983 -1165 4075 -1159
rect 3983 -1199 3995 -1165
rect 4063 -1199 4075 -1165
rect 3983 -1205 4075 -1199
rect 4141 -1165 4233 -1159
rect 4141 -1199 4153 -1165
rect 4221 -1199 4233 -1165
rect 4141 -1205 4233 -1199
rect 4299 -1165 4391 -1159
rect 4299 -1199 4311 -1165
rect 4379 -1199 4391 -1165
rect 4299 -1205 4391 -1199
rect 4457 -1165 4549 -1159
rect 4457 -1199 4469 -1165
rect 4537 -1199 4549 -1165
rect 4457 -1205 4549 -1199
rect 4615 -1165 4707 -1159
rect 4615 -1199 4627 -1165
rect 4695 -1199 4707 -1165
rect 4615 -1205 4707 -1199
rect 4773 -1165 4865 -1159
rect 4773 -1199 4785 -1165
rect 4853 -1199 4865 -1165
rect 4773 -1205 4865 -1199
rect -4865 -1273 -4773 -1267
rect -4865 -1307 -4853 -1273
rect -4785 -1307 -4773 -1273
rect -4865 -1313 -4773 -1307
rect -4707 -1273 -4615 -1267
rect -4707 -1307 -4695 -1273
rect -4627 -1307 -4615 -1273
rect -4707 -1313 -4615 -1307
rect -4549 -1273 -4457 -1267
rect -4549 -1307 -4537 -1273
rect -4469 -1307 -4457 -1273
rect -4549 -1313 -4457 -1307
rect -4391 -1273 -4299 -1267
rect -4391 -1307 -4379 -1273
rect -4311 -1307 -4299 -1273
rect -4391 -1313 -4299 -1307
rect -4233 -1273 -4141 -1267
rect -4233 -1307 -4221 -1273
rect -4153 -1307 -4141 -1273
rect -4233 -1313 -4141 -1307
rect -4075 -1273 -3983 -1267
rect -4075 -1307 -4063 -1273
rect -3995 -1307 -3983 -1273
rect -4075 -1313 -3983 -1307
rect -3917 -1273 -3825 -1267
rect -3917 -1307 -3905 -1273
rect -3837 -1307 -3825 -1273
rect -3917 -1313 -3825 -1307
rect -3759 -1273 -3667 -1267
rect -3759 -1307 -3747 -1273
rect -3679 -1307 -3667 -1273
rect -3759 -1313 -3667 -1307
rect -3601 -1273 -3509 -1267
rect -3601 -1307 -3589 -1273
rect -3521 -1307 -3509 -1273
rect -3601 -1313 -3509 -1307
rect -3443 -1273 -3351 -1267
rect -3443 -1307 -3431 -1273
rect -3363 -1307 -3351 -1273
rect -3443 -1313 -3351 -1307
rect -3285 -1273 -3193 -1267
rect -3285 -1307 -3273 -1273
rect -3205 -1307 -3193 -1273
rect -3285 -1313 -3193 -1307
rect -3127 -1273 -3035 -1267
rect -3127 -1307 -3115 -1273
rect -3047 -1307 -3035 -1273
rect -3127 -1313 -3035 -1307
rect -2969 -1273 -2877 -1267
rect -2969 -1307 -2957 -1273
rect -2889 -1307 -2877 -1273
rect -2969 -1313 -2877 -1307
rect -2811 -1273 -2719 -1267
rect -2811 -1307 -2799 -1273
rect -2731 -1307 -2719 -1273
rect -2811 -1313 -2719 -1307
rect -2653 -1273 -2561 -1267
rect -2653 -1307 -2641 -1273
rect -2573 -1307 -2561 -1273
rect -2653 -1313 -2561 -1307
rect -2495 -1273 -2403 -1267
rect -2495 -1307 -2483 -1273
rect -2415 -1307 -2403 -1273
rect -2495 -1313 -2403 -1307
rect -2337 -1273 -2245 -1267
rect -2337 -1307 -2325 -1273
rect -2257 -1307 -2245 -1273
rect -2337 -1313 -2245 -1307
rect -2179 -1273 -2087 -1267
rect -2179 -1307 -2167 -1273
rect -2099 -1307 -2087 -1273
rect -2179 -1313 -2087 -1307
rect -2021 -1273 -1929 -1267
rect -2021 -1307 -2009 -1273
rect -1941 -1307 -1929 -1273
rect -2021 -1313 -1929 -1307
rect -1863 -1273 -1771 -1267
rect -1863 -1307 -1851 -1273
rect -1783 -1307 -1771 -1273
rect -1863 -1313 -1771 -1307
rect -1705 -1273 -1613 -1267
rect -1705 -1307 -1693 -1273
rect -1625 -1307 -1613 -1273
rect -1705 -1313 -1613 -1307
rect -1547 -1273 -1455 -1267
rect -1547 -1307 -1535 -1273
rect -1467 -1307 -1455 -1273
rect -1547 -1313 -1455 -1307
rect -1389 -1273 -1297 -1267
rect -1389 -1307 -1377 -1273
rect -1309 -1307 -1297 -1273
rect -1389 -1313 -1297 -1307
rect -1231 -1273 -1139 -1267
rect -1231 -1307 -1219 -1273
rect -1151 -1307 -1139 -1273
rect -1231 -1313 -1139 -1307
rect -1073 -1273 -981 -1267
rect -1073 -1307 -1061 -1273
rect -993 -1307 -981 -1273
rect -1073 -1313 -981 -1307
rect -915 -1273 -823 -1267
rect -915 -1307 -903 -1273
rect -835 -1307 -823 -1273
rect -915 -1313 -823 -1307
rect -757 -1273 -665 -1267
rect -757 -1307 -745 -1273
rect -677 -1307 -665 -1273
rect -757 -1313 -665 -1307
rect -599 -1273 -507 -1267
rect -599 -1307 -587 -1273
rect -519 -1307 -507 -1273
rect -599 -1313 -507 -1307
rect -441 -1273 -349 -1267
rect -441 -1307 -429 -1273
rect -361 -1307 -349 -1273
rect -441 -1313 -349 -1307
rect -283 -1273 -191 -1267
rect -283 -1307 -271 -1273
rect -203 -1307 -191 -1273
rect -283 -1313 -191 -1307
rect -125 -1273 -33 -1267
rect -125 -1307 -113 -1273
rect -45 -1307 -33 -1273
rect -125 -1313 -33 -1307
rect 33 -1273 125 -1267
rect 33 -1307 45 -1273
rect 113 -1307 125 -1273
rect 33 -1313 125 -1307
rect 191 -1273 283 -1267
rect 191 -1307 203 -1273
rect 271 -1307 283 -1273
rect 191 -1313 283 -1307
rect 349 -1273 441 -1267
rect 349 -1307 361 -1273
rect 429 -1307 441 -1273
rect 349 -1313 441 -1307
rect 507 -1273 599 -1267
rect 507 -1307 519 -1273
rect 587 -1307 599 -1273
rect 507 -1313 599 -1307
rect 665 -1273 757 -1267
rect 665 -1307 677 -1273
rect 745 -1307 757 -1273
rect 665 -1313 757 -1307
rect 823 -1273 915 -1267
rect 823 -1307 835 -1273
rect 903 -1307 915 -1273
rect 823 -1313 915 -1307
rect 981 -1273 1073 -1267
rect 981 -1307 993 -1273
rect 1061 -1307 1073 -1273
rect 981 -1313 1073 -1307
rect 1139 -1273 1231 -1267
rect 1139 -1307 1151 -1273
rect 1219 -1307 1231 -1273
rect 1139 -1313 1231 -1307
rect 1297 -1273 1389 -1267
rect 1297 -1307 1309 -1273
rect 1377 -1307 1389 -1273
rect 1297 -1313 1389 -1307
rect 1455 -1273 1547 -1267
rect 1455 -1307 1467 -1273
rect 1535 -1307 1547 -1273
rect 1455 -1313 1547 -1307
rect 1613 -1273 1705 -1267
rect 1613 -1307 1625 -1273
rect 1693 -1307 1705 -1273
rect 1613 -1313 1705 -1307
rect 1771 -1273 1863 -1267
rect 1771 -1307 1783 -1273
rect 1851 -1307 1863 -1273
rect 1771 -1313 1863 -1307
rect 1929 -1273 2021 -1267
rect 1929 -1307 1941 -1273
rect 2009 -1307 2021 -1273
rect 1929 -1313 2021 -1307
rect 2087 -1273 2179 -1267
rect 2087 -1307 2099 -1273
rect 2167 -1307 2179 -1273
rect 2087 -1313 2179 -1307
rect 2245 -1273 2337 -1267
rect 2245 -1307 2257 -1273
rect 2325 -1307 2337 -1273
rect 2245 -1313 2337 -1307
rect 2403 -1273 2495 -1267
rect 2403 -1307 2415 -1273
rect 2483 -1307 2495 -1273
rect 2403 -1313 2495 -1307
rect 2561 -1273 2653 -1267
rect 2561 -1307 2573 -1273
rect 2641 -1307 2653 -1273
rect 2561 -1313 2653 -1307
rect 2719 -1273 2811 -1267
rect 2719 -1307 2731 -1273
rect 2799 -1307 2811 -1273
rect 2719 -1313 2811 -1307
rect 2877 -1273 2969 -1267
rect 2877 -1307 2889 -1273
rect 2957 -1307 2969 -1273
rect 2877 -1313 2969 -1307
rect 3035 -1273 3127 -1267
rect 3035 -1307 3047 -1273
rect 3115 -1307 3127 -1273
rect 3035 -1313 3127 -1307
rect 3193 -1273 3285 -1267
rect 3193 -1307 3205 -1273
rect 3273 -1307 3285 -1273
rect 3193 -1313 3285 -1307
rect 3351 -1273 3443 -1267
rect 3351 -1307 3363 -1273
rect 3431 -1307 3443 -1273
rect 3351 -1313 3443 -1307
rect 3509 -1273 3601 -1267
rect 3509 -1307 3521 -1273
rect 3589 -1307 3601 -1273
rect 3509 -1313 3601 -1307
rect 3667 -1273 3759 -1267
rect 3667 -1307 3679 -1273
rect 3747 -1307 3759 -1273
rect 3667 -1313 3759 -1307
rect 3825 -1273 3917 -1267
rect 3825 -1307 3837 -1273
rect 3905 -1307 3917 -1273
rect 3825 -1313 3917 -1307
rect 3983 -1273 4075 -1267
rect 3983 -1307 3995 -1273
rect 4063 -1307 4075 -1273
rect 3983 -1313 4075 -1307
rect 4141 -1273 4233 -1267
rect 4141 -1307 4153 -1273
rect 4221 -1307 4233 -1273
rect 4141 -1313 4233 -1307
rect 4299 -1273 4391 -1267
rect 4299 -1307 4311 -1273
rect 4379 -1307 4391 -1273
rect 4299 -1313 4391 -1307
rect 4457 -1273 4549 -1267
rect 4457 -1307 4469 -1273
rect 4537 -1307 4549 -1273
rect 4457 -1313 4549 -1307
rect 4615 -1273 4707 -1267
rect 4615 -1307 4627 -1273
rect 4695 -1307 4707 -1273
rect 4615 -1313 4707 -1307
rect 4773 -1273 4865 -1267
rect 4773 -1307 4785 -1273
rect 4853 -1307 4865 -1273
rect 4773 -1313 4865 -1307
rect -4921 -1366 -4875 -1354
rect -4921 -2342 -4915 -1366
rect -4881 -2342 -4875 -1366
rect -4921 -2354 -4875 -2342
rect -4763 -1366 -4717 -1354
rect -4763 -2342 -4757 -1366
rect -4723 -2342 -4717 -1366
rect -4763 -2354 -4717 -2342
rect -4605 -1366 -4559 -1354
rect -4605 -2342 -4599 -1366
rect -4565 -2342 -4559 -1366
rect -4605 -2354 -4559 -2342
rect -4447 -1366 -4401 -1354
rect -4447 -2342 -4441 -1366
rect -4407 -2342 -4401 -1366
rect -4447 -2354 -4401 -2342
rect -4289 -1366 -4243 -1354
rect -4289 -2342 -4283 -1366
rect -4249 -2342 -4243 -1366
rect -4289 -2354 -4243 -2342
rect -4131 -1366 -4085 -1354
rect -4131 -2342 -4125 -1366
rect -4091 -2342 -4085 -1366
rect -4131 -2354 -4085 -2342
rect -3973 -1366 -3927 -1354
rect -3973 -2342 -3967 -1366
rect -3933 -2342 -3927 -1366
rect -3973 -2354 -3927 -2342
rect -3815 -1366 -3769 -1354
rect -3815 -2342 -3809 -1366
rect -3775 -2342 -3769 -1366
rect -3815 -2354 -3769 -2342
rect -3657 -1366 -3611 -1354
rect -3657 -2342 -3651 -1366
rect -3617 -2342 -3611 -1366
rect -3657 -2354 -3611 -2342
rect -3499 -1366 -3453 -1354
rect -3499 -2342 -3493 -1366
rect -3459 -2342 -3453 -1366
rect -3499 -2354 -3453 -2342
rect -3341 -1366 -3295 -1354
rect -3341 -2342 -3335 -1366
rect -3301 -2342 -3295 -1366
rect -3341 -2354 -3295 -2342
rect -3183 -1366 -3137 -1354
rect -3183 -2342 -3177 -1366
rect -3143 -2342 -3137 -1366
rect -3183 -2354 -3137 -2342
rect -3025 -1366 -2979 -1354
rect -3025 -2342 -3019 -1366
rect -2985 -2342 -2979 -1366
rect -3025 -2354 -2979 -2342
rect -2867 -1366 -2821 -1354
rect -2867 -2342 -2861 -1366
rect -2827 -2342 -2821 -1366
rect -2867 -2354 -2821 -2342
rect -2709 -1366 -2663 -1354
rect -2709 -2342 -2703 -1366
rect -2669 -2342 -2663 -1366
rect -2709 -2354 -2663 -2342
rect -2551 -1366 -2505 -1354
rect -2551 -2342 -2545 -1366
rect -2511 -2342 -2505 -1366
rect -2551 -2354 -2505 -2342
rect -2393 -1366 -2347 -1354
rect -2393 -2342 -2387 -1366
rect -2353 -2342 -2347 -1366
rect -2393 -2354 -2347 -2342
rect -2235 -1366 -2189 -1354
rect -2235 -2342 -2229 -1366
rect -2195 -2342 -2189 -1366
rect -2235 -2354 -2189 -2342
rect -2077 -1366 -2031 -1354
rect -2077 -2342 -2071 -1366
rect -2037 -2342 -2031 -1366
rect -2077 -2354 -2031 -2342
rect -1919 -1366 -1873 -1354
rect -1919 -2342 -1913 -1366
rect -1879 -2342 -1873 -1366
rect -1919 -2354 -1873 -2342
rect -1761 -1366 -1715 -1354
rect -1761 -2342 -1755 -1366
rect -1721 -2342 -1715 -1366
rect -1761 -2354 -1715 -2342
rect -1603 -1366 -1557 -1354
rect -1603 -2342 -1597 -1366
rect -1563 -2342 -1557 -1366
rect -1603 -2354 -1557 -2342
rect -1445 -1366 -1399 -1354
rect -1445 -2342 -1439 -1366
rect -1405 -2342 -1399 -1366
rect -1445 -2354 -1399 -2342
rect -1287 -1366 -1241 -1354
rect -1287 -2342 -1281 -1366
rect -1247 -2342 -1241 -1366
rect -1287 -2354 -1241 -2342
rect -1129 -1366 -1083 -1354
rect -1129 -2342 -1123 -1366
rect -1089 -2342 -1083 -1366
rect -1129 -2354 -1083 -2342
rect -971 -1366 -925 -1354
rect -971 -2342 -965 -1366
rect -931 -2342 -925 -1366
rect -971 -2354 -925 -2342
rect -813 -1366 -767 -1354
rect -813 -2342 -807 -1366
rect -773 -2342 -767 -1366
rect -813 -2354 -767 -2342
rect -655 -1366 -609 -1354
rect -655 -2342 -649 -1366
rect -615 -2342 -609 -1366
rect -655 -2354 -609 -2342
rect -497 -1366 -451 -1354
rect -497 -2342 -491 -1366
rect -457 -2342 -451 -1366
rect -497 -2354 -451 -2342
rect -339 -1366 -293 -1354
rect -339 -2342 -333 -1366
rect -299 -2342 -293 -1366
rect -339 -2354 -293 -2342
rect -181 -1366 -135 -1354
rect -181 -2342 -175 -1366
rect -141 -2342 -135 -1366
rect -181 -2354 -135 -2342
rect -23 -1366 23 -1354
rect -23 -2342 -17 -1366
rect 17 -2342 23 -1366
rect -23 -2354 23 -2342
rect 135 -1366 181 -1354
rect 135 -2342 141 -1366
rect 175 -2342 181 -1366
rect 135 -2354 181 -2342
rect 293 -1366 339 -1354
rect 293 -2342 299 -1366
rect 333 -2342 339 -1366
rect 293 -2354 339 -2342
rect 451 -1366 497 -1354
rect 451 -2342 457 -1366
rect 491 -2342 497 -1366
rect 451 -2354 497 -2342
rect 609 -1366 655 -1354
rect 609 -2342 615 -1366
rect 649 -2342 655 -1366
rect 609 -2354 655 -2342
rect 767 -1366 813 -1354
rect 767 -2342 773 -1366
rect 807 -2342 813 -1366
rect 767 -2354 813 -2342
rect 925 -1366 971 -1354
rect 925 -2342 931 -1366
rect 965 -2342 971 -1366
rect 925 -2354 971 -2342
rect 1083 -1366 1129 -1354
rect 1083 -2342 1089 -1366
rect 1123 -2342 1129 -1366
rect 1083 -2354 1129 -2342
rect 1241 -1366 1287 -1354
rect 1241 -2342 1247 -1366
rect 1281 -2342 1287 -1366
rect 1241 -2354 1287 -2342
rect 1399 -1366 1445 -1354
rect 1399 -2342 1405 -1366
rect 1439 -2342 1445 -1366
rect 1399 -2354 1445 -2342
rect 1557 -1366 1603 -1354
rect 1557 -2342 1563 -1366
rect 1597 -2342 1603 -1366
rect 1557 -2354 1603 -2342
rect 1715 -1366 1761 -1354
rect 1715 -2342 1721 -1366
rect 1755 -2342 1761 -1366
rect 1715 -2354 1761 -2342
rect 1873 -1366 1919 -1354
rect 1873 -2342 1879 -1366
rect 1913 -2342 1919 -1366
rect 1873 -2354 1919 -2342
rect 2031 -1366 2077 -1354
rect 2031 -2342 2037 -1366
rect 2071 -2342 2077 -1366
rect 2031 -2354 2077 -2342
rect 2189 -1366 2235 -1354
rect 2189 -2342 2195 -1366
rect 2229 -2342 2235 -1366
rect 2189 -2354 2235 -2342
rect 2347 -1366 2393 -1354
rect 2347 -2342 2353 -1366
rect 2387 -2342 2393 -1366
rect 2347 -2354 2393 -2342
rect 2505 -1366 2551 -1354
rect 2505 -2342 2511 -1366
rect 2545 -2342 2551 -1366
rect 2505 -2354 2551 -2342
rect 2663 -1366 2709 -1354
rect 2663 -2342 2669 -1366
rect 2703 -2342 2709 -1366
rect 2663 -2354 2709 -2342
rect 2821 -1366 2867 -1354
rect 2821 -2342 2827 -1366
rect 2861 -2342 2867 -1366
rect 2821 -2354 2867 -2342
rect 2979 -1366 3025 -1354
rect 2979 -2342 2985 -1366
rect 3019 -2342 3025 -1366
rect 2979 -2354 3025 -2342
rect 3137 -1366 3183 -1354
rect 3137 -2342 3143 -1366
rect 3177 -2342 3183 -1366
rect 3137 -2354 3183 -2342
rect 3295 -1366 3341 -1354
rect 3295 -2342 3301 -1366
rect 3335 -2342 3341 -1366
rect 3295 -2354 3341 -2342
rect 3453 -1366 3499 -1354
rect 3453 -2342 3459 -1366
rect 3493 -2342 3499 -1366
rect 3453 -2354 3499 -2342
rect 3611 -1366 3657 -1354
rect 3611 -2342 3617 -1366
rect 3651 -2342 3657 -1366
rect 3611 -2354 3657 -2342
rect 3769 -1366 3815 -1354
rect 3769 -2342 3775 -1366
rect 3809 -2342 3815 -1366
rect 3769 -2354 3815 -2342
rect 3927 -1366 3973 -1354
rect 3927 -2342 3933 -1366
rect 3967 -2342 3973 -1366
rect 3927 -2354 3973 -2342
rect 4085 -1366 4131 -1354
rect 4085 -2342 4091 -1366
rect 4125 -2342 4131 -1366
rect 4085 -2354 4131 -2342
rect 4243 -1366 4289 -1354
rect 4243 -2342 4249 -1366
rect 4283 -2342 4289 -1366
rect 4243 -2354 4289 -2342
rect 4401 -1366 4447 -1354
rect 4401 -2342 4407 -1366
rect 4441 -2342 4447 -1366
rect 4401 -2354 4447 -2342
rect 4559 -1366 4605 -1354
rect 4559 -2342 4565 -1366
rect 4599 -2342 4605 -1366
rect 4559 -2354 4605 -2342
rect 4717 -1366 4763 -1354
rect 4717 -2342 4723 -1366
rect 4757 -2342 4763 -1366
rect 4717 -2354 4763 -2342
rect 4875 -1366 4921 -1354
rect 4875 -2342 4881 -1366
rect 4915 -2342 4921 -1366
rect 4875 -2354 4921 -2342
rect -4865 -2401 -4773 -2395
rect -4865 -2435 -4853 -2401
rect -4785 -2435 -4773 -2401
rect -4865 -2441 -4773 -2435
rect -4707 -2401 -4615 -2395
rect -4707 -2435 -4695 -2401
rect -4627 -2435 -4615 -2401
rect -4707 -2441 -4615 -2435
rect -4549 -2401 -4457 -2395
rect -4549 -2435 -4537 -2401
rect -4469 -2435 -4457 -2401
rect -4549 -2441 -4457 -2435
rect -4391 -2401 -4299 -2395
rect -4391 -2435 -4379 -2401
rect -4311 -2435 -4299 -2401
rect -4391 -2441 -4299 -2435
rect -4233 -2401 -4141 -2395
rect -4233 -2435 -4221 -2401
rect -4153 -2435 -4141 -2401
rect -4233 -2441 -4141 -2435
rect -4075 -2401 -3983 -2395
rect -4075 -2435 -4063 -2401
rect -3995 -2435 -3983 -2401
rect -4075 -2441 -3983 -2435
rect -3917 -2401 -3825 -2395
rect -3917 -2435 -3905 -2401
rect -3837 -2435 -3825 -2401
rect -3917 -2441 -3825 -2435
rect -3759 -2401 -3667 -2395
rect -3759 -2435 -3747 -2401
rect -3679 -2435 -3667 -2401
rect -3759 -2441 -3667 -2435
rect -3601 -2401 -3509 -2395
rect -3601 -2435 -3589 -2401
rect -3521 -2435 -3509 -2401
rect -3601 -2441 -3509 -2435
rect -3443 -2401 -3351 -2395
rect -3443 -2435 -3431 -2401
rect -3363 -2435 -3351 -2401
rect -3443 -2441 -3351 -2435
rect -3285 -2401 -3193 -2395
rect -3285 -2435 -3273 -2401
rect -3205 -2435 -3193 -2401
rect -3285 -2441 -3193 -2435
rect -3127 -2401 -3035 -2395
rect -3127 -2435 -3115 -2401
rect -3047 -2435 -3035 -2401
rect -3127 -2441 -3035 -2435
rect -2969 -2401 -2877 -2395
rect -2969 -2435 -2957 -2401
rect -2889 -2435 -2877 -2401
rect -2969 -2441 -2877 -2435
rect -2811 -2401 -2719 -2395
rect -2811 -2435 -2799 -2401
rect -2731 -2435 -2719 -2401
rect -2811 -2441 -2719 -2435
rect -2653 -2401 -2561 -2395
rect -2653 -2435 -2641 -2401
rect -2573 -2435 -2561 -2401
rect -2653 -2441 -2561 -2435
rect -2495 -2401 -2403 -2395
rect -2495 -2435 -2483 -2401
rect -2415 -2435 -2403 -2401
rect -2495 -2441 -2403 -2435
rect -2337 -2401 -2245 -2395
rect -2337 -2435 -2325 -2401
rect -2257 -2435 -2245 -2401
rect -2337 -2441 -2245 -2435
rect -2179 -2401 -2087 -2395
rect -2179 -2435 -2167 -2401
rect -2099 -2435 -2087 -2401
rect -2179 -2441 -2087 -2435
rect -2021 -2401 -1929 -2395
rect -2021 -2435 -2009 -2401
rect -1941 -2435 -1929 -2401
rect -2021 -2441 -1929 -2435
rect -1863 -2401 -1771 -2395
rect -1863 -2435 -1851 -2401
rect -1783 -2435 -1771 -2401
rect -1863 -2441 -1771 -2435
rect -1705 -2401 -1613 -2395
rect -1705 -2435 -1693 -2401
rect -1625 -2435 -1613 -2401
rect -1705 -2441 -1613 -2435
rect -1547 -2401 -1455 -2395
rect -1547 -2435 -1535 -2401
rect -1467 -2435 -1455 -2401
rect -1547 -2441 -1455 -2435
rect -1389 -2401 -1297 -2395
rect -1389 -2435 -1377 -2401
rect -1309 -2435 -1297 -2401
rect -1389 -2441 -1297 -2435
rect -1231 -2401 -1139 -2395
rect -1231 -2435 -1219 -2401
rect -1151 -2435 -1139 -2401
rect -1231 -2441 -1139 -2435
rect -1073 -2401 -981 -2395
rect -1073 -2435 -1061 -2401
rect -993 -2435 -981 -2401
rect -1073 -2441 -981 -2435
rect -915 -2401 -823 -2395
rect -915 -2435 -903 -2401
rect -835 -2435 -823 -2401
rect -915 -2441 -823 -2435
rect -757 -2401 -665 -2395
rect -757 -2435 -745 -2401
rect -677 -2435 -665 -2401
rect -757 -2441 -665 -2435
rect -599 -2401 -507 -2395
rect -599 -2435 -587 -2401
rect -519 -2435 -507 -2401
rect -599 -2441 -507 -2435
rect -441 -2401 -349 -2395
rect -441 -2435 -429 -2401
rect -361 -2435 -349 -2401
rect -441 -2441 -349 -2435
rect -283 -2401 -191 -2395
rect -283 -2435 -271 -2401
rect -203 -2435 -191 -2401
rect -283 -2441 -191 -2435
rect -125 -2401 -33 -2395
rect -125 -2435 -113 -2401
rect -45 -2435 -33 -2401
rect -125 -2441 -33 -2435
rect 33 -2401 125 -2395
rect 33 -2435 45 -2401
rect 113 -2435 125 -2401
rect 33 -2441 125 -2435
rect 191 -2401 283 -2395
rect 191 -2435 203 -2401
rect 271 -2435 283 -2401
rect 191 -2441 283 -2435
rect 349 -2401 441 -2395
rect 349 -2435 361 -2401
rect 429 -2435 441 -2401
rect 349 -2441 441 -2435
rect 507 -2401 599 -2395
rect 507 -2435 519 -2401
rect 587 -2435 599 -2401
rect 507 -2441 599 -2435
rect 665 -2401 757 -2395
rect 665 -2435 677 -2401
rect 745 -2435 757 -2401
rect 665 -2441 757 -2435
rect 823 -2401 915 -2395
rect 823 -2435 835 -2401
rect 903 -2435 915 -2401
rect 823 -2441 915 -2435
rect 981 -2401 1073 -2395
rect 981 -2435 993 -2401
rect 1061 -2435 1073 -2401
rect 981 -2441 1073 -2435
rect 1139 -2401 1231 -2395
rect 1139 -2435 1151 -2401
rect 1219 -2435 1231 -2401
rect 1139 -2441 1231 -2435
rect 1297 -2401 1389 -2395
rect 1297 -2435 1309 -2401
rect 1377 -2435 1389 -2401
rect 1297 -2441 1389 -2435
rect 1455 -2401 1547 -2395
rect 1455 -2435 1467 -2401
rect 1535 -2435 1547 -2401
rect 1455 -2441 1547 -2435
rect 1613 -2401 1705 -2395
rect 1613 -2435 1625 -2401
rect 1693 -2435 1705 -2401
rect 1613 -2441 1705 -2435
rect 1771 -2401 1863 -2395
rect 1771 -2435 1783 -2401
rect 1851 -2435 1863 -2401
rect 1771 -2441 1863 -2435
rect 1929 -2401 2021 -2395
rect 1929 -2435 1941 -2401
rect 2009 -2435 2021 -2401
rect 1929 -2441 2021 -2435
rect 2087 -2401 2179 -2395
rect 2087 -2435 2099 -2401
rect 2167 -2435 2179 -2401
rect 2087 -2441 2179 -2435
rect 2245 -2401 2337 -2395
rect 2245 -2435 2257 -2401
rect 2325 -2435 2337 -2401
rect 2245 -2441 2337 -2435
rect 2403 -2401 2495 -2395
rect 2403 -2435 2415 -2401
rect 2483 -2435 2495 -2401
rect 2403 -2441 2495 -2435
rect 2561 -2401 2653 -2395
rect 2561 -2435 2573 -2401
rect 2641 -2435 2653 -2401
rect 2561 -2441 2653 -2435
rect 2719 -2401 2811 -2395
rect 2719 -2435 2731 -2401
rect 2799 -2435 2811 -2401
rect 2719 -2441 2811 -2435
rect 2877 -2401 2969 -2395
rect 2877 -2435 2889 -2401
rect 2957 -2435 2969 -2401
rect 2877 -2441 2969 -2435
rect 3035 -2401 3127 -2395
rect 3035 -2435 3047 -2401
rect 3115 -2435 3127 -2401
rect 3035 -2441 3127 -2435
rect 3193 -2401 3285 -2395
rect 3193 -2435 3205 -2401
rect 3273 -2435 3285 -2401
rect 3193 -2441 3285 -2435
rect 3351 -2401 3443 -2395
rect 3351 -2435 3363 -2401
rect 3431 -2435 3443 -2401
rect 3351 -2441 3443 -2435
rect 3509 -2401 3601 -2395
rect 3509 -2435 3521 -2401
rect 3589 -2435 3601 -2401
rect 3509 -2441 3601 -2435
rect 3667 -2401 3759 -2395
rect 3667 -2435 3679 -2401
rect 3747 -2435 3759 -2401
rect 3667 -2441 3759 -2435
rect 3825 -2401 3917 -2395
rect 3825 -2435 3837 -2401
rect 3905 -2435 3917 -2401
rect 3825 -2441 3917 -2435
rect 3983 -2401 4075 -2395
rect 3983 -2435 3995 -2401
rect 4063 -2435 4075 -2401
rect 3983 -2441 4075 -2435
rect 4141 -2401 4233 -2395
rect 4141 -2435 4153 -2401
rect 4221 -2435 4233 -2401
rect 4141 -2441 4233 -2435
rect 4299 -2401 4391 -2395
rect 4299 -2435 4311 -2401
rect 4379 -2435 4391 -2401
rect 4299 -2441 4391 -2435
rect 4457 -2401 4549 -2395
rect 4457 -2435 4469 -2401
rect 4537 -2435 4549 -2401
rect 4457 -2441 4549 -2435
rect 4615 -2401 4707 -2395
rect 4615 -2435 4627 -2401
rect 4695 -2435 4707 -2401
rect 4615 -2441 4707 -2435
rect 4773 -2401 4865 -2395
rect 4773 -2435 4785 -2401
rect 4853 -2435 4865 -2401
rect 4773 -2441 4865 -2435
<< properties >>
string FIXED_BBOX -5032 -2556 5032 2556
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.5 m 4 nf 62 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
