magic
tech sky130A
magscale 1 2
timestamp 1757105855
<< nwell >>
rect -3583 -797 3583 797
<< mvpmos >>
rect -3325 -500 -3125 500
rect -3067 -500 -2867 500
rect -2809 -500 -2609 500
rect -2551 -500 -2351 500
rect -2293 -500 -2093 500
rect -2035 -500 -1835 500
rect -1777 -500 -1577 500
rect -1519 -500 -1319 500
rect -1261 -500 -1061 500
rect -1003 -500 -803 500
rect -745 -500 -545 500
rect -487 -500 -287 500
rect -229 -500 -29 500
rect 29 -500 229 500
rect 287 -500 487 500
rect 545 -500 745 500
rect 803 -500 1003 500
rect 1061 -500 1261 500
rect 1319 -500 1519 500
rect 1577 -500 1777 500
rect 1835 -500 2035 500
rect 2093 -500 2293 500
rect 2351 -500 2551 500
rect 2609 -500 2809 500
rect 2867 -500 3067 500
rect 3125 -500 3325 500
<< mvpdiff >>
rect -3383 488 -3325 500
rect -3383 -488 -3371 488
rect -3337 -488 -3325 488
rect -3383 -500 -3325 -488
rect -3125 488 -3067 500
rect -3125 -488 -3113 488
rect -3079 -488 -3067 488
rect -3125 -500 -3067 -488
rect -2867 488 -2809 500
rect -2867 -488 -2855 488
rect -2821 -488 -2809 488
rect -2867 -500 -2809 -488
rect -2609 488 -2551 500
rect -2609 -488 -2597 488
rect -2563 -488 -2551 488
rect -2609 -500 -2551 -488
rect -2351 488 -2293 500
rect -2351 -488 -2339 488
rect -2305 -488 -2293 488
rect -2351 -500 -2293 -488
rect -2093 488 -2035 500
rect -2093 -488 -2081 488
rect -2047 -488 -2035 488
rect -2093 -500 -2035 -488
rect -1835 488 -1777 500
rect -1835 -488 -1823 488
rect -1789 -488 -1777 488
rect -1835 -500 -1777 -488
rect -1577 488 -1519 500
rect -1577 -488 -1565 488
rect -1531 -488 -1519 488
rect -1577 -500 -1519 -488
rect -1319 488 -1261 500
rect -1319 -488 -1307 488
rect -1273 -488 -1261 488
rect -1319 -500 -1261 -488
rect -1061 488 -1003 500
rect -1061 -488 -1049 488
rect -1015 -488 -1003 488
rect -1061 -500 -1003 -488
rect -803 488 -745 500
rect -803 -488 -791 488
rect -757 -488 -745 488
rect -803 -500 -745 -488
rect -545 488 -487 500
rect -545 -488 -533 488
rect -499 -488 -487 488
rect -545 -500 -487 -488
rect -287 488 -229 500
rect -287 -488 -275 488
rect -241 -488 -229 488
rect -287 -500 -229 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 229 488 287 500
rect 229 -488 241 488
rect 275 -488 287 488
rect 229 -500 287 -488
rect 487 488 545 500
rect 487 -488 499 488
rect 533 -488 545 488
rect 487 -500 545 -488
rect 745 488 803 500
rect 745 -488 757 488
rect 791 -488 803 488
rect 745 -500 803 -488
rect 1003 488 1061 500
rect 1003 -488 1015 488
rect 1049 -488 1061 488
rect 1003 -500 1061 -488
rect 1261 488 1319 500
rect 1261 -488 1273 488
rect 1307 -488 1319 488
rect 1261 -500 1319 -488
rect 1519 488 1577 500
rect 1519 -488 1531 488
rect 1565 -488 1577 488
rect 1519 -500 1577 -488
rect 1777 488 1835 500
rect 1777 -488 1789 488
rect 1823 -488 1835 488
rect 1777 -500 1835 -488
rect 2035 488 2093 500
rect 2035 -488 2047 488
rect 2081 -488 2093 488
rect 2035 -500 2093 -488
rect 2293 488 2351 500
rect 2293 -488 2305 488
rect 2339 -488 2351 488
rect 2293 -500 2351 -488
rect 2551 488 2609 500
rect 2551 -488 2563 488
rect 2597 -488 2609 488
rect 2551 -500 2609 -488
rect 2809 488 2867 500
rect 2809 -488 2821 488
rect 2855 -488 2867 488
rect 2809 -500 2867 -488
rect 3067 488 3125 500
rect 3067 -488 3079 488
rect 3113 -488 3125 488
rect 3067 -500 3125 -488
rect 3325 488 3383 500
rect 3325 -488 3337 488
rect 3371 -488 3383 488
rect 3325 -500 3383 -488
<< mvpdiffc >>
rect -3371 -488 -3337 488
rect -3113 -488 -3079 488
rect -2855 -488 -2821 488
rect -2597 -488 -2563 488
rect -2339 -488 -2305 488
rect -2081 -488 -2047 488
rect -1823 -488 -1789 488
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect 1789 -488 1823 488
rect 2047 -488 2081 488
rect 2305 -488 2339 488
rect 2563 -488 2597 488
rect 2821 -488 2855 488
rect 3079 -488 3113 488
rect 3337 -488 3371 488
<< mvnsubdiff >>
rect -3517 719 3517 731
rect -3517 685 -3409 719
rect 3409 685 3517 719
rect -3517 673 3517 685
rect -3517 623 -3459 673
rect -3517 -623 -3505 623
rect -3471 -623 -3459 623
rect 3459 623 3517 673
rect -3517 -673 -3459 -623
rect 3459 -623 3471 623
rect 3505 -623 3517 623
rect 3459 -673 3517 -623
rect -3517 -685 3517 -673
rect -3517 -719 -3409 -685
rect 3409 -719 3517 -685
rect -3517 -731 3517 -719
<< mvnsubdiffcont >>
rect -3409 685 3409 719
rect -3505 -623 -3471 623
rect 3471 -623 3505 623
rect -3409 -719 3409 -685
<< poly >>
rect -3325 581 -3125 597
rect -3325 547 -3309 581
rect -3141 547 -3125 581
rect -3325 500 -3125 547
rect -3067 581 -2867 597
rect -3067 547 -3051 581
rect -2883 547 -2867 581
rect -3067 500 -2867 547
rect -2809 581 -2609 597
rect -2809 547 -2793 581
rect -2625 547 -2609 581
rect -2809 500 -2609 547
rect -2551 581 -2351 597
rect -2551 547 -2535 581
rect -2367 547 -2351 581
rect -2551 500 -2351 547
rect -2293 581 -2093 597
rect -2293 547 -2277 581
rect -2109 547 -2093 581
rect -2293 500 -2093 547
rect -2035 581 -1835 597
rect -2035 547 -2019 581
rect -1851 547 -1835 581
rect -2035 500 -1835 547
rect -1777 581 -1577 597
rect -1777 547 -1761 581
rect -1593 547 -1577 581
rect -1777 500 -1577 547
rect -1519 581 -1319 597
rect -1519 547 -1503 581
rect -1335 547 -1319 581
rect -1519 500 -1319 547
rect -1261 581 -1061 597
rect -1261 547 -1245 581
rect -1077 547 -1061 581
rect -1261 500 -1061 547
rect -1003 581 -803 597
rect -1003 547 -987 581
rect -819 547 -803 581
rect -1003 500 -803 547
rect -745 581 -545 597
rect -745 547 -729 581
rect -561 547 -545 581
rect -745 500 -545 547
rect -487 581 -287 597
rect -487 547 -471 581
rect -303 547 -287 581
rect -487 500 -287 547
rect -229 581 -29 597
rect -229 547 -213 581
rect -45 547 -29 581
rect -229 500 -29 547
rect 29 581 229 597
rect 29 547 45 581
rect 213 547 229 581
rect 29 500 229 547
rect 287 581 487 597
rect 287 547 303 581
rect 471 547 487 581
rect 287 500 487 547
rect 545 581 745 597
rect 545 547 561 581
rect 729 547 745 581
rect 545 500 745 547
rect 803 581 1003 597
rect 803 547 819 581
rect 987 547 1003 581
rect 803 500 1003 547
rect 1061 581 1261 597
rect 1061 547 1077 581
rect 1245 547 1261 581
rect 1061 500 1261 547
rect 1319 581 1519 597
rect 1319 547 1335 581
rect 1503 547 1519 581
rect 1319 500 1519 547
rect 1577 581 1777 597
rect 1577 547 1593 581
rect 1761 547 1777 581
rect 1577 500 1777 547
rect 1835 581 2035 597
rect 1835 547 1851 581
rect 2019 547 2035 581
rect 1835 500 2035 547
rect 2093 581 2293 597
rect 2093 547 2109 581
rect 2277 547 2293 581
rect 2093 500 2293 547
rect 2351 581 2551 597
rect 2351 547 2367 581
rect 2535 547 2551 581
rect 2351 500 2551 547
rect 2609 581 2809 597
rect 2609 547 2625 581
rect 2793 547 2809 581
rect 2609 500 2809 547
rect 2867 581 3067 597
rect 2867 547 2883 581
rect 3051 547 3067 581
rect 2867 500 3067 547
rect 3125 581 3325 597
rect 3125 547 3141 581
rect 3309 547 3325 581
rect 3125 500 3325 547
rect -3325 -547 -3125 -500
rect -3325 -581 -3309 -547
rect -3141 -581 -3125 -547
rect -3325 -597 -3125 -581
rect -3067 -547 -2867 -500
rect -3067 -581 -3051 -547
rect -2883 -581 -2867 -547
rect -3067 -597 -2867 -581
rect -2809 -547 -2609 -500
rect -2809 -581 -2793 -547
rect -2625 -581 -2609 -547
rect -2809 -597 -2609 -581
rect -2551 -547 -2351 -500
rect -2551 -581 -2535 -547
rect -2367 -581 -2351 -547
rect -2551 -597 -2351 -581
rect -2293 -547 -2093 -500
rect -2293 -581 -2277 -547
rect -2109 -581 -2093 -547
rect -2293 -597 -2093 -581
rect -2035 -547 -1835 -500
rect -2035 -581 -2019 -547
rect -1851 -581 -1835 -547
rect -2035 -597 -1835 -581
rect -1777 -547 -1577 -500
rect -1777 -581 -1761 -547
rect -1593 -581 -1577 -547
rect -1777 -597 -1577 -581
rect -1519 -547 -1319 -500
rect -1519 -581 -1503 -547
rect -1335 -581 -1319 -547
rect -1519 -597 -1319 -581
rect -1261 -547 -1061 -500
rect -1261 -581 -1245 -547
rect -1077 -581 -1061 -547
rect -1261 -597 -1061 -581
rect -1003 -547 -803 -500
rect -1003 -581 -987 -547
rect -819 -581 -803 -547
rect -1003 -597 -803 -581
rect -745 -547 -545 -500
rect -745 -581 -729 -547
rect -561 -581 -545 -547
rect -745 -597 -545 -581
rect -487 -547 -287 -500
rect -487 -581 -471 -547
rect -303 -581 -287 -547
rect -487 -597 -287 -581
rect -229 -547 -29 -500
rect -229 -581 -213 -547
rect -45 -581 -29 -547
rect -229 -597 -29 -581
rect 29 -547 229 -500
rect 29 -581 45 -547
rect 213 -581 229 -547
rect 29 -597 229 -581
rect 287 -547 487 -500
rect 287 -581 303 -547
rect 471 -581 487 -547
rect 287 -597 487 -581
rect 545 -547 745 -500
rect 545 -581 561 -547
rect 729 -581 745 -547
rect 545 -597 745 -581
rect 803 -547 1003 -500
rect 803 -581 819 -547
rect 987 -581 1003 -547
rect 803 -597 1003 -581
rect 1061 -547 1261 -500
rect 1061 -581 1077 -547
rect 1245 -581 1261 -547
rect 1061 -597 1261 -581
rect 1319 -547 1519 -500
rect 1319 -581 1335 -547
rect 1503 -581 1519 -547
rect 1319 -597 1519 -581
rect 1577 -547 1777 -500
rect 1577 -581 1593 -547
rect 1761 -581 1777 -547
rect 1577 -597 1777 -581
rect 1835 -547 2035 -500
rect 1835 -581 1851 -547
rect 2019 -581 2035 -547
rect 1835 -597 2035 -581
rect 2093 -547 2293 -500
rect 2093 -581 2109 -547
rect 2277 -581 2293 -547
rect 2093 -597 2293 -581
rect 2351 -547 2551 -500
rect 2351 -581 2367 -547
rect 2535 -581 2551 -547
rect 2351 -597 2551 -581
rect 2609 -547 2809 -500
rect 2609 -581 2625 -547
rect 2793 -581 2809 -547
rect 2609 -597 2809 -581
rect 2867 -547 3067 -500
rect 2867 -581 2883 -547
rect 3051 -581 3067 -547
rect 2867 -597 3067 -581
rect 3125 -547 3325 -500
rect 3125 -581 3141 -547
rect 3309 -581 3325 -547
rect 3125 -597 3325 -581
<< polycont >>
rect -3309 547 -3141 581
rect -3051 547 -2883 581
rect -2793 547 -2625 581
rect -2535 547 -2367 581
rect -2277 547 -2109 581
rect -2019 547 -1851 581
rect -1761 547 -1593 581
rect -1503 547 -1335 581
rect -1245 547 -1077 581
rect -987 547 -819 581
rect -729 547 -561 581
rect -471 547 -303 581
rect -213 547 -45 581
rect 45 547 213 581
rect 303 547 471 581
rect 561 547 729 581
rect 819 547 987 581
rect 1077 547 1245 581
rect 1335 547 1503 581
rect 1593 547 1761 581
rect 1851 547 2019 581
rect 2109 547 2277 581
rect 2367 547 2535 581
rect 2625 547 2793 581
rect 2883 547 3051 581
rect 3141 547 3309 581
rect -3309 -581 -3141 -547
rect -3051 -581 -2883 -547
rect -2793 -581 -2625 -547
rect -2535 -581 -2367 -547
rect -2277 -581 -2109 -547
rect -2019 -581 -1851 -547
rect -1761 -581 -1593 -547
rect -1503 -581 -1335 -547
rect -1245 -581 -1077 -547
rect -987 -581 -819 -547
rect -729 -581 -561 -547
rect -471 -581 -303 -547
rect -213 -581 -45 -547
rect 45 -581 213 -547
rect 303 -581 471 -547
rect 561 -581 729 -547
rect 819 -581 987 -547
rect 1077 -581 1245 -547
rect 1335 -581 1503 -547
rect 1593 -581 1761 -547
rect 1851 -581 2019 -547
rect 2109 -581 2277 -547
rect 2367 -581 2535 -547
rect 2625 -581 2793 -547
rect 2883 -581 3051 -547
rect 3141 -581 3309 -547
<< locali >>
rect -3505 685 -3409 719
rect 3409 685 3505 719
rect -3505 623 -3471 685
rect 3471 623 3505 685
rect -3325 547 -3309 581
rect -3141 547 -3125 581
rect -3067 547 -3051 581
rect -2883 547 -2867 581
rect -2809 547 -2793 581
rect -2625 547 -2609 581
rect -2551 547 -2535 581
rect -2367 547 -2351 581
rect -2293 547 -2277 581
rect -2109 547 -2093 581
rect -2035 547 -2019 581
rect -1851 547 -1835 581
rect -1777 547 -1761 581
rect -1593 547 -1577 581
rect -1519 547 -1503 581
rect -1335 547 -1319 581
rect -1261 547 -1245 581
rect -1077 547 -1061 581
rect -1003 547 -987 581
rect -819 547 -803 581
rect -745 547 -729 581
rect -561 547 -545 581
rect -487 547 -471 581
rect -303 547 -287 581
rect -229 547 -213 581
rect -45 547 -29 581
rect 29 547 45 581
rect 213 547 229 581
rect 287 547 303 581
rect 471 547 487 581
rect 545 547 561 581
rect 729 547 745 581
rect 803 547 819 581
rect 987 547 1003 581
rect 1061 547 1077 581
rect 1245 547 1261 581
rect 1319 547 1335 581
rect 1503 547 1519 581
rect 1577 547 1593 581
rect 1761 547 1777 581
rect 1835 547 1851 581
rect 2019 547 2035 581
rect 2093 547 2109 581
rect 2277 547 2293 581
rect 2351 547 2367 581
rect 2535 547 2551 581
rect 2609 547 2625 581
rect 2793 547 2809 581
rect 2867 547 2883 581
rect 3051 547 3067 581
rect 3125 547 3141 581
rect 3309 547 3325 581
rect -3371 488 -3337 504
rect -3371 -504 -3337 -488
rect -3113 488 -3079 504
rect -3113 -504 -3079 -488
rect -2855 488 -2821 504
rect -2855 -504 -2821 -488
rect -2597 488 -2563 504
rect -2597 -504 -2563 -488
rect -2339 488 -2305 504
rect -2339 -504 -2305 -488
rect -2081 488 -2047 504
rect -2081 -504 -2047 -488
rect -1823 488 -1789 504
rect -1823 -504 -1789 -488
rect -1565 488 -1531 504
rect -1565 -504 -1531 -488
rect -1307 488 -1273 504
rect -1307 -504 -1273 -488
rect -1049 488 -1015 504
rect -1049 -504 -1015 -488
rect -791 488 -757 504
rect -791 -504 -757 -488
rect -533 488 -499 504
rect -533 -504 -499 -488
rect -275 488 -241 504
rect -275 -504 -241 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 241 488 275 504
rect 241 -504 275 -488
rect 499 488 533 504
rect 499 -504 533 -488
rect 757 488 791 504
rect 757 -504 791 -488
rect 1015 488 1049 504
rect 1015 -504 1049 -488
rect 1273 488 1307 504
rect 1273 -504 1307 -488
rect 1531 488 1565 504
rect 1531 -504 1565 -488
rect 1789 488 1823 504
rect 1789 -504 1823 -488
rect 2047 488 2081 504
rect 2047 -504 2081 -488
rect 2305 488 2339 504
rect 2305 -504 2339 -488
rect 2563 488 2597 504
rect 2563 -504 2597 -488
rect 2821 488 2855 504
rect 2821 -504 2855 -488
rect 3079 488 3113 504
rect 3079 -504 3113 -488
rect 3337 488 3371 504
rect 3337 -504 3371 -488
rect -3325 -581 -3309 -547
rect -3141 -581 -3125 -547
rect -3067 -581 -3051 -547
rect -2883 -581 -2867 -547
rect -2809 -581 -2793 -547
rect -2625 -581 -2609 -547
rect -2551 -581 -2535 -547
rect -2367 -581 -2351 -547
rect -2293 -581 -2277 -547
rect -2109 -581 -2093 -547
rect -2035 -581 -2019 -547
rect -1851 -581 -1835 -547
rect -1777 -581 -1761 -547
rect -1593 -581 -1577 -547
rect -1519 -581 -1503 -547
rect -1335 -581 -1319 -547
rect -1261 -581 -1245 -547
rect -1077 -581 -1061 -547
rect -1003 -581 -987 -547
rect -819 -581 -803 -547
rect -745 -581 -729 -547
rect -561 -581 -545 -547
rect -487 -581 -471 -547
rect -303 -581 -287 -547
rect -229 -581 -213 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 213 -581 229 -547
rect 287 -581 303 -547
rect 471 -581 487 -547
rect 545 -581 561 -547
rect 729 -581 745 -547
rect 803 -581 819 -547
rect 987 -581 1003 -547
rect 1061 -581 1077 -547
rect 1245 -581 1261 -547
rect 1319 -581 1335 -547
rect 1503 -581 1519 -547
rect 1577 -581 1593 -547
rect 1761 -581 1777 -547
rect 1835 -581 1851 -547
rect 2019 -581 2035 -547
rect 2093 -581 2109 -547
rect 2277 -581 2293 -547
rect 2351 -581 2367 -547
rect 2535 -581 2551 -547
rect 2609 -581 2625 -547
rect 2793 -581 2809 -547
rect 2867 -581 2883 -547
rect 3051 -581 3067 -547
rect 3125 -581 3141 -547
rect 3309 -581 3325 -547
rect -3505 -685 -3471 -623
rect 3471 -685 3505 -623
rect -3505 -719 -3409 -685
rect 3409 -719 3505 -685
<< viali >>
rect -3309 547 -3141 581
rect -3051 547 -2883 581
rect -2793 547 -2625 581
rect -2535 547 -2367 581
rect -2277 547 -2109 581
rect -2019 547 -1851 581
rect -1761 547 -1593 581
rect -1503 547 -1335 581
rect -1245 547 -1077 581
rect -987 547 -819 581
rect -729 547 -561 581
rect -471 547 -303 581
rect -213 547 -45 581
rect 45 547 213 581
rect 303 547 471 581
rect 561 547 729 581
rect 819 547 987 581
rect 1077 547 1245 581
rect 1335 547 1503 581
rect 1593 547 1761 581
rect 1851 547 2019 581
rect 2109 547 2277 581
rect 2367 547 2535 581
rect 2625 547 2793 581
rect 2883 547 3051 581
rect 3141 547 3309 581
rect -3371 -488 -3337 488
rect -3113 -488 -3079 488
rect -2855 -488 -2821 488
rect -2597 -488 -2563 488
rect -2339 -488 -2305 488
rect -2081 -488 -2047 488
rect -1823 -488 -1789 488
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect 1789 -488 1823 488
rect 2047 -488 2081 488
rect 2305 -488 2339 488
rect 2563 -488 2597 488
rect 2821 -488 2855 488
rect 3079 -488 3113 488
rect 3337 -488 3371 488
rect -3309 -581 -3141 -547
rect -3051 -581 -2883 -547
rect -2793 -581 -2625 -547
rect -2535 -581 -2367 -547
rect -2277 -581 -2109 -547
rect -2019 -581 -1851 -547
rect -1761 -581 -1593 -547
rect -1503 -581 -1335 -547
rect -1245 -581 -1077 -547
rect -987 -581 -819 -547
rect -729 -581 -561 -547
rect -471 -581 -303 -547
rect -213 -581 -45 -547
rect 45 -581 213 -547
rect 303 -581 471 -547
rect 561 -581 729 -547
rect 819 -581 987 -547
rect 1077 -581 1245 -547
rect 1335 -581 1503 -547
rect 1593 -581 1761 -547
rect 1851 -581 2019 -547
rect 2109 -581 2277 -547
rect 2367 -581 2535 -547
rect 2625 -581 2793 -547
rect 2883 -581 3051 -547
rect 3141 -581 3309 -547
<< metal1 >>
rect -3321 581 -3129 587
rect -3321 547 -3309 581
rect -3141 547 -3129 581
rect -3321 541 -3129 547
rect -3063 581 -2871 587
rect -3063 547 -3051 581
rect -2883 547 -2871 581
rect -3063 541 -2871 547
rect -2805 581 -2613 587
rect -2805 547 -2793 581
rect -2625 547 -2613 581
rect -2805 541 -2613 547
rect -2547 581 -2355 587
rect -2547 547 -2535 581
rect -2367 547 -2355 581
rect -2547 541 -2355 547
rect -2289 581 -2097 587
rect -2289 547 -2277 581
rect -2109 547 -2097 581
rect -2289 541 -2097 547
rect -2031 581 -1839 587
rect -2031 547 -2019 581
rect -1851 547 -1839 581
rect -2031 541 -1839 547
rect -1773 581 -1581 587
rect -1773 547 -1761 581
rect -1593 547 -1581 581
rect -1773 541 -1581 547
rect -1515 581 -1323 587
rect -1515 547 -1503 581
rect -1335 547 -1323 581
rect -1515 541 -1323 547
rect -1257 581 -1065 587
rect -1257 547 -1245 581
rect -1077 547 -1065 581
rect -1257 541 -1065 547
rect -999 581 -807 587
rect -999 547 -987 581
rect -819 547 -807 581
rect -999 541 -807 547
rect -741 581 -549 587
rect -741 547 -729 581
rect -561 547 -549 581
rect -741 541 -549 547
rect -483 581 -291 587
rect -483 547 -471 581
rect -303 547 -291 581
rect -483 541 -291 547
rect -225 581 -33 587
rect -225 547 -213 581
rect -45 547 -33 581
rect -225 541 -33 547
rect 33 581 225 587
rect 33 547 45 581
rect 213 547 225 581
rect 33 541 225 547
rect 291 581 483 587
rect 291 547 303 581
rect 471 547 483 581
rect 291 541 483 547
rect 549 581 741 587
rect 549 547 561 581
rect 729 547 741 581
rect 549 541 741 547
rect 807 581 999 587
rect 807 547 819 581
rect 987 547 999 581
rect 807 541 999 547
rect 1065 581 1257 587
rect 1065 547 1077 581
rect 1245 547 1257 581
rect 1065 541 1257 547
rect 1323 581 1515 587
rect 1323 547 1335 581
rect 1503 547 1515 581
rect 1323 541 1515 547
rect 1581 581 1773 587
rect 1581 547 1593 581
rect 1761 547 1773 581
rect 1581 541 1773 547
rect 1839 581 2031 587
rect 1839 547 1851 581
rect 2019 547 2031 581
rect 1839 541 2031 547
rect 2097 581 2289 587
rect 2097 547 2109 581
rect 2277 547 2289 581
rect 2097 541 2289 547
rect 2355 581 2547 587
rect 2355 547 2367 581
rect 2535 547 2547 581
rect 2355 541 2547 547
rect 2613 581 2805 587
rect 2613 547 2625 581
rect 2793 547 2805 581
rect 2613 541 2805 547
rect 2871 581 3063 587
rect 2871 547 2883 581
rect 3051 547 3063 581
rect 2871 541 3063 547
rect 3129 581 3321 587
rect 3129 547 3141 581
rect 3309 547 3321 581
rect 3129 541 3321 547
rect -3377 488 -3331 500
rect -3377 -488 -3371 488
rect -3337 -488 -3331 488
rect -3377 -500 -3331 -488
rect -3119 488 -3073 500
rect -3119 -488 -3113 488
rect -3079 -488 -3073 488
rect -3119 -500 -3073 -488
rect -2861 488 -2815 500
rect -2861 -488 -2855 488
rect -2821 -488 -2815 488
rect -2861 -500 -2815 -488
rect -2603 488 -2557 500
rect -2603 -488 -2597 488
rect -2563 -488 -2557 488
rect -2603 -500 -2557 -488
rect -2345 488 -2299 500
rect -2345 -488 -2339 488
rect -2305 -488 -2299 488
rect -2345 -500 -2299 -488
rect -2087 488 -2041 500
rect -2087 -488 -2081 488
rect -2047 -488 -2041 488
rect -2087 -500 -2041 -488
rect -1829 488 -1783 500
rect -1829 -488 -1823 488
rect -1789 -488 -1783 488
rect -1829 -500 -1783 -488
rect -1571 488 -1525 500
rect -1571 -488 -1565 488
rect -1531 -488 -1525 488
rect -1571 -500 -1525 -488
rect -1313 488 -1267 500
rect -1313 -488 -1307 488
rect -1273 -488 -1267 488
rect -1313 -500 -1267 -488
rect -1055 488 -1009 500
rect -1055 -488 -1049 488
rect -1015 -488 -1009 488
rect -1055 -500 -1009 -488
rect -797 488 -751 500
rect -797 -488 -791 488
rect -757 -488 -751 488
rect -797 -500 -751 -488
rect -539 488 -493 500
rect -539 -488 -533 488
rect -499 -488 -493 488
rect -539 -500 -493 -488
rect -281 488 -235 500
rect -281 -488 -275 488
rect -241 -488 -235 488
rect -281 -500 -235 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 235 488 281 500
rect 235 -488 241 488
rect 275 -488 281 488
rect 235 -500 281 -488
rect 493 488 539 500
rect 493 -488 499 488
rect 533 -488 539 488
rect 493 -500 539 -488
rect 751 488 797 500
rect 751 -488 757 488
rect 791 -488 797 488
rect 751 -500 797 -488
rect 1009 488 1055 500
rect 1009 -488 1015 488
rect 1049 -488 1055 488
rect 1009 -500 1055 -488
rect 1267 488 1313 500
rect 1267 -488 1273 488
rect 1307 -488 1313 488
rect 1267 -500 1313 -488
rect 1525 488 1571 500
rect 1525 -488 1531 488
rect 1565 -488 1571 488
rect 1525 -500 1571 -488
rect 1783 488 1829 500
rect 1783 -488 1789 488
rect 1823 -488 1829 488
rect 1783 -500 1829 -488
rect 2041 488 2087 500
rect 2041 -488 2047 488
rect 2081 -488 2087 488
rect 2041 -500 2087 -488
rect 2299 488 2345 500
rect 2299 -488 2305 488
rect 2339 -488 2345 488
rect 2299 -500 2345 -488
rect 2557 488 2603 500
rect 2557 -488 2563 488
rect 2597 -488 2603 488
rect 2557 -500 2603 -488
rect 2815 488 2861 500
rect 2815 -488 2821 488
rect 2855 -488 2861 488
rect 2815 -500 2861 -488
rect 3073 488 3119 500
rect 3073 -488 3079 488
rect 3113 -488 3119 488
rect 3073 -500 3119 -488
rect 3331 488 3377 500
rect 3331 -488 3337 488
rect 3371 -488 3377 488
rect 3331 -500 3377 -488
rect -3321 -547 -3129 -541
rect -3321 -581 -3309 -547
rect -3141 -581 -3129 -547
rect -3321 -587 -3129 -581
rect -3063 -547 -2871 -541
rect -3063 -581 -3051 -547
rect -2883 -581 -2871 -547
rect -3063 -587 -2871 -581
rect -2805 -547 -2613 -541
rect -2805 -581 -2793 -547
rect -2625 -581 -2613 -547
rect -2805 -587 -2613 -581
rect -2547 -547 -2355 -541
rect -2547 -581 -2535 -547
rect -2367 -581 -2355 -547
rect -2547 -587 -2355 -581
rect -2289 -547 -2097 -541
rect -2289 -581 -2277 -547
rect -2109 -581 -2097 -547
rect -2289 -587 -2097 -581
rect -2031 -547 -1839 -541
rect -2031 -581 -2019 -547
rect -1851 -581 -1839 -547
rect -2031 -587 -1839 -581
rect -1773 -547 -1581 -541
rect -1773 -581 -1761 -547
rect -1593 -581 -1581 -547
rect -1773 -587 -1581 -581
rect -1515 -547 -1323 -541
rect -1515 -581 -1503 -547
rect -1335 -581 -1323 -547
rect -1515 -587 -1323 -581
rect -1257 -547 -1065 -541
rect -1257 -581 -1245 -547
rect -1077 -581 -1065 -547
rect -1257 -587 -1065 -581
rect -999 -547 -807 -541
rect -999 -581 -987 -547
rect -819 -581 -807 -547
rect -999 -587 -807 -581
rect -741 -547 -549 -541
rect -741 -581 -729 -547
rect -561 -581 -549 -547
rect -741 -587 -549 -581
rect -483 -547 -291 -541
rect -483 -581 -471 -547
rect -303 -581 -291 -547
rect -483 -587 -291 -581
rect -225 -547 -33 -541
rect -225 -581 -213 -547
rect -45 -581 -33 -547
rect -225 -587 -33 -581
rect 33 -547 225 -541
rect 33 -581 45 -547
rect 213 -581 225 -547
rect 33 -587 225 -581
rect 291 -547 483 -541
rect 291 -581 303 -547
rect 471 -581 483 -547
rect 291 -587 483 -581
rect 549 -547 741 -541
rect 549 -581 561 -547
rect 729 -581 741 -547
rect 549 -587 741 -581
rect 807 -547 999 -541
rect 807 -581 819 -547
rect 987 -581 999 -547
rect 807 -587 999 -581
rect 1065 -547 1257 -541
rect 1065 -581 1077 -547
rect 1245 -581 1257 -547
rect 1065 -587 1257 -581
rect 1323 -547 1515 -541
rect 1323 -581 1335 -547
rect 1503 -581 1515 -547
rect 1323 -587 1515 -581
rect 1581 -547 1773 -541
rect 1581 -581 1593 -547
rect 1761 -581 1773 -547
rect 1581 -587 1773 -581
rect 1839 -547 2031 -541
rect 1839 -581 1851 -547
rect 2019 -581 2031 -547
rect 1839 -587 2031 -581
rect 2097 -547 2289 -541
rect 2097 -581 2109 -547
rect 2277 -581 2289 -547
rect 2097 -587 2289 -581
rect 2355 -547 2547 -541
rect 2355 -581 2367 -547
rect 2535 -581 2547 -547
rect 2355 -587 2547 -581
rect 2613 -547 2805 -541
rect 2613 -581 2625 -547
rect 2793 -581 2805 -547
rect 2613 -587 2805 -581
rect 2871 -547 3063 -541
rect 2871 -581 2883 -547
rect 3051 -581 3063 -547
rect 2871 -587 3063 -581
rect 3129 -547 3321 -541
rect 3129 -581 3141 -547
rect 3309 -581 3321 -547
rect 3129 -587 3321 -581
<< properties >>
string FIXED_BBOX -3488 -702 3488 702
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 1 m 1 nf 26 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
