** sch_path: /foss/designs/ttsky25a_minimosbius/xschem/tb_mosbius_dpn_dc.sch
**.subckt tb_mosbius_dpn_dc
x1 g g g g g g VAPWR v g g v g g VDPWR GND net1[4] net1[3] net1[2] net1[1] net1[0] v g g v g g g g g
+ v g g g g g v g g g g g v g g GND GND GND g g g v g g g g g v g g g g v g v g g g v g g g net2 g v g
+ g g g GND GND GND GND GND GND GND GND v g g v g g g g g v g g g g g v g g g g g v g g g g g v g g g g
+ g v g g GND GND vs1 vs0 g g g v g g GND GND g g g v g g g g g v g g g g g v g g g g g v g g g g g v g
+ g GND GND g g g v g g GND GND GND GND g g g v g g g g g v g g GND GND GND GND GND GND v v v v v v v v
+ v v v mosbius
VAPWR VAPWR GND 3.3
.save i(vapwr)
VDPWR VDPWR GND 1.8
.save i(vdpwr)
Ibias GND Ibias 100u
VSIG vsig GND 0
.save i(vsig)
VCM net3 GND 1.8
.save i(vcm)
R13 g GND 1u m=1
R14 v VDPWR 1u m=1
x3 VAPWR VDPWR ibias_ref GND GND GND GND GND GND GND GND mirror_n
Ibias1 GND ibias_ref 100u
x2[5] GND voutm net1[4] pad_model
x2[4] GND voutp net1[3] pad_model
x2[3] GND g net1[2] pad_model
x2[2] GND vinm net1[1] pad_model
x2[1] GND vinp net1[0] pad_model
x2 GND Ibias net2 pad_model
Vmeasm VAPWR voutm 0
.save i(vmeasm)
Vmeasp VAPWR voutp 0
.save i(vmeasp)
x4 VAPWR VDPWR net4 net5 vinp vinm vs1 vs0 GND ibias_ref GND diff_n
Vmeasp_ref VAPWR net4 0
.save i(vmeasp_ref)
Vmeasm_ref VAPWR net5 0
.save i(vmeasm_ref)
E1 vinm net3 vsig GND -0.5
E2 vinp net3 vsig GND 0.5
VS1 vs1 GND 0
.save i(vs1)
VS0 vs0 GND 0
.save i(vs0)
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice



*****************************************
* MOSBIUS: N-Diff Pair DC Test
*****************************************
* output current vs input voltage for the n-chnl differential pair.
* compares the dp with mosbius parasitics vs dp in isolation
* steps through tail current values.
* plots iout vs vin and gm vs vin
*****************************************
* BUS1: DP INP
* BUS2: DP INM
* BUS3: GND
* BUS4: DP OUTP
* BUS5: DP OUTM
* BUS6: GND
*****************************************
.control
   save all
   set temp = 27
   repeat 2
      repeat 2
         dc vsig -1 1 0.01
         alter VS0 1.8
      end
      alter VS0 0
      alter VS1 1.8
   end
   let mosb_200u = dc1.i(vmeasp)-dc1.i(vmeasm)
   let base_200u = dc1.i(vmeasp_ref)-dc1.i(vmeasm_ref)
   let mosb_400u = dc2.i(vmeasp)-dc2.i(vmeasm)
   let base_400u = dc2.i(vmeasp_ref)-dc2.i(vmeasm_ref)
   let mosb_600u = dc3.i(vmeasp)-dc3.i(vmeasm)
   let base_600u = dc3.i(vmeasp_ref)-dc3.i(vmeasm_ref)
   let mosb_800u = dc4.i(vmeasp)-dc4.i(vmeasm)
   let base_800u = dc4.i(vmeasp_ref)-dc4.i(vmeasm_ref)
   let mosb_gm_200u = deriv(mosb_200u)
   let base_gm_200u = deriv(base_200u)
   let mosb_gm_400u = deriv(mosb_400u)
   let base_gm_400u = deriv(base_400u)
   let mosb_gm_600u = deriv(mosb_600u)
   let base_gm_600u = deriv(base_600u)
   let mosb_gm_800u = deriv(mosb_800u)
   let base_gm_800u = deriv(base_800u)
   plot mosb_200u base_200u mosb_400u base_400u mosb_600u base_600u mosb_800u base_800u
   plot mosb_gm_200u base_gm_200u mosb_gm_400u base_gm_400u mosb_gm_600u base_gm_600u mosb_gm_800u
+ base_gm_800u
.endc


**** end user architecture code
**.ends

* expanding   symbol:  mosbius.sym # of pins=54
** sym_path: /foss/designs/ttsky25a_minimosbius/xschem/mosbius.sym
** sch_path: /foss/designs/ttsky25a_minimosbius/xschem/mosbius.sch
.subckt mosbius cfga_vapwr[6] cfga_vapwr[5] cfga_vapwr[4] cfga_vapwr[3] cfga_vapwr[2] cfga_vapwr[1]
+ VAPWR cfga_vgnd[6] cfga_vgnd[5] cfga_vgnd[4] cfga_vgnd[3] cfga_vgnd[2] cfga_vgnd[1] VDPWR VGND bus_A[5]
+ bus_A[4] bus_A[3] bus_A[2] bus_A[1] cfga_otan_inp[3] cfga_otan_inp[2] cfga_otan_inp[1] cfgb_otan_inm[3]
+ cfgb_otan_inm[2] cfgb_otan_inm[1] cfga_otan_out[6] cfga_otan_out[5] cfga_otan_out[4] cfga_otan_out[3]
+ cfga_otan_out[2] cfga_otan_out[1] cfga_mirn_a[6] cfga_mirn_a[5] cfga_mirn_a[4] cfga_mirn_a[3] cfga_mirn_a[2]
+ cfga_mirn_a[1] cfgb_mirn_b[6] cfgb_mirn_b[5] cfgb_mirn_b[4] cfgb_mirn_b[3] cfgb_mirn_b[2] cfgb_mirn_b[1]
+ ctrl_otan_tail[1] ctrl_otan_tail[0] ctrl_otan_diode cfga_mirp_a[6] cfga_mirp_a[5] cfga_mirp_a[4] cfga_mirp_a[3]
+ cfga_mirp_a[2] cfga_mirp_a[1] cfgb_mirp_b[6] cfgb_mirp_b[5] cfgb_mirp_b[4] cfgb_mirp_b[3] cfgb_mirp_b[2]
+ cfgb_mirp_b[1] cfga_dpn_inp[3] cfga_dpn_inp[2] cfga_dpn_inp[1] cfgb_dpn_inm[3] cfgb_dpn_inm[2] cfgb_dpn_inm[1]
+ cfga_dpn_outp[6] cfga_dpn_outp[5] cfga_dpn_outp[4] cfga_dpn_outp[3] cfga_dpn_outp[2] cfga_dpn_outp[1] ibias
+ cfgb_dpn_outm[6] cfgb_dpn_outm[5] cfgb_dpn_outm[4] cfgb_dpn_outm[3] cfgb_dpn_outm[2] cfgb_dpn_outm[1] ctrl_mirp_a[1]
+ ctrl_mirp_a[0] ctrl_mirn_a[1] ctrl_mirn_a[0] ctrl_mirp_b[1] ctrl_mirp_b[0] ctrl_mirn_b[1] ctrl_mirn_b[0]
+ cfga_dpp_inp[3] cfga_dpp_inp[2] cfga_dpp_inp[1] cfgb_dpp_inm[3] cfgb_dpp_inm[2] cfgb_dpp_inm[1] cfga_dpp_outp[6]
+ cfga_dpp_outp[5] cfga_dpp_outp[4] cfga_dpp_outp[3] cfga_dpp_outp[2] cfga_dpp_outp[1] cfgb_dpp_outm[6]
+ cfgb_dpp_outm[5] cfgb_dpp_outm[4] cfgb_dpp_outm[3] cfgb_dpp_outm[2] cfgb_dpp_outm[1] cfga_nfeta_d[6] cfga_nfeta_d[5]
+ cfga_nfeta_d[4] cfga_nfeta_d[3] cfga_nfeta_d[2] cfga_nfeta_d[1] cfgb_nfetb_d[6] cfgb_nfetb_d[5] cfgb_nfetb_d[4]
+ cfgb_nfetb_d[3] cfgb_nfetb_d[2] cfgb_nfetb_d[1] cfga_nfeta_g[6] cfga_nfeta_g[5] cfga_nfeta_g[4] cfga_nfeta_g[3]
+ cfga_nfeta_g[2] cfga_nfeta_g[1] ctrl_dpp_tail[1] ctrl_dpp_tail[0] ctrl_dpn_tail[1] ctrl_dpn_tail[0] cfgb_nfetb_g[6]
+ cfgb_nfetb_g[5] cfgb_nfetb_g[4] cfgb_nfetb_g[3] cfgb_nfetb_g[2] cfgb_nfetb_g[1] ctrl_dpp_source ctrl_dpn_source
+ cfga_nfeta_s[6] cfga_nfeta_s[5] cfga_nfeta_s[4] cfga_nfeta_s[3] cfga_nfeta_s[2] cfga_nfeta_s[1] cfgb_nfetb_s[6]
+ cfgb_nfetb_s[5] cfgb_nfetb_s[4] cfgb_nfetb_s[3] cfgb_nfetb_s[2] cfgb_nfetb_s[1] cfga_pfeta_d[6] cfga_pfeta_d[5]
+ cfga_pfeta_d[4] cfga_pfeta_d[3] cfga_pfeta_d[2] cfga_pfeta_d[1] cfgb_pfetb_d[6] cfgb_pfetb_d[5] cfgb_pfetb_d[4]
+ cfgb_pfetb_d[3] cfgb_pfetb_d[2] cfgb_pfetb_d[1] cfga_pfeta_g[6] cfga_pfeta_g[5] cfga_pfeta_g[4] cfga_pfeta_g[3]
+ cfga_pfeta_g[2] cfga_pfeta_g[1] ctrl_pfeta_source ctrl_nfeta_source cfgb_pfetb_g[6] cfgb_pfetb_g[5] cfgb_pfetb_g[4]
+ cfgb_pfetb_g[3] cfgb_pfetb_g[2] cfgb_pfetb_g[1] ctrl_pfeta_width[1] ctrl_pfeta_width[0] ctrl_nfeta_width[1]
+ ctrl_nfeta_width[0] cfga_pfeta_s[6] cfga_pfeta_s[5] cfga_pfeta_s[4] cfga_pfeta_s[3] cfga_pfeta_s[2] cfga_pfeta_s[1]
+ cfgb_pfetb_s[6] cfgb_pfetb_s[5] cfgb_pfetb_s[4] cfgb_pfetb_s[3] cfgb_pfetb_s[2] cfgb_pfetb_s[1] ctrl_pfetb_source
+ ctrl_nfetb_source ctrl_pfetb_width[1] ctrl_pfetb_width[0] ctrl_nfetb_width[1] ctrl_nfetb_width[0] cfg_bus_short[6]
+ cfg_bus_short[5] cfg_bus_short[4] cfg_bus_short[3] cfg_bus_short[2] cfg_bus_short[1] cfg_bus_ext[5] cfg_bus_ext[4]
+ cfg_bus_ext[3] cfg_bus_ext[2] cfg_bus_ext[1]
*.ipin cfga_vapwr[6],cfga_vapwr[5],cfga_vapwr[4],cfga_vapwr[3],cfga_vapwr[2],cfga_vapwr[1]
*.ipin cfga_vgnd[6],cfga_vgnd[5],cfga_vgnd[4],cfga_vgnd[3],cfga_vgnd[2],cfga_vgnd[1]
*.ipin cfga_otan_inp[3],cfga_otan_inp[2],cfga_otan_inp[1]
*.ipin
*+ cfga_otan_out[6],cfga_otan_out[5],cfga_otan_out[4],cfga_otan_out[3],cfga_otan_out[2],cfga_otan_out[1]
*.ipin cfga_mirn_a[6],cfga_mirn_a[5],cfga_mirn_a[4],cfga_mirn_a[3],cfga_mirn_a[2],cfga_mirn_a[1]
*.ipin cfga_mirp_a[6],cfga_mirp_a[5],cfga_mirp_a[4],cfga_mirp_a[3],cfga_mirp_a[2],cfga_mirp_a[1]
*.ipin cfga_dpn_inp[3],cfga_dpn_inp[2],cfga_dpn_inp[1]
*.ipin
*+ cfga_dpn_outp[6],cfga_dpn_outp[5],cfga_dpn_outp[4],cfga_dpn_outp[3],cfga_dpn_outp[2],cfga_dpn_outp[1]
*.ipin cfga_dpp_inp[3],cfga_dpp_inp[2],cfga_dpp_inp[1]
*.ipin
*+ cfga_dpp_outp[6],cfga_dpp_outp[5],cfga_dpp_outp[4],cfga_dpp_outp[3],cfga_dpp_outp[2],cfga_dpp_outp[1]
*.ipin
*+ cfga_nfeta_d[6],cfga_nfeta_d[5],cfga_nfeta_d[4],cfga_nfeta_d[3],cfga_nfeta_d[2],cfga_nfeta_d[1]
*.ipin
*+ cfga_nfeta_g[6],cfga_nfeta_g[5],cfga_nfeta_g[4],cfga_nfeta_g[3],cfga_nfeta_g[2],cfga_nfeta_g[1]
*.ipin
*+ cfga_nfeta_s[6],cfga_nfeta_s[5],cfga_nfeta_s[4],cfga_nfeta_s[3],cfga_nfeta_s[2],cfga_nfeta_s[1]
*.ipin
*+ cfga_pfeta_d[6],cfga_pfeta_d[5],cfga_pfeta_d[4],cfga_pfeta_d[3],cfga_pfeta_d[2],cfga_pfeta_d[1]
*.ipin
*+ cfga_pfeta_g[6],cfga_pfeta_g[5],cfga_pfeta_g[4],cfga_pfeta_g[3],cfga_pfeta_g[2],cfga_pfeta_g[1]
*.ipin
*+ cfga_pfeta_s[6],cfga_pfeta_s[5],cfga_pfeta_s[4],cfga_pfeta_s[3],cfga_pfeta_s[2],cfga_pfeta_s[1]
*.ipin cfgb_otan_inm[3],cfgb_otan_inm[2],cfgb_otan_inm[1]
*.ipin cfgb_mirn_b[6],cfgb_mirn_b[5],cfgb_mirn_b[4],cfgb_mirn_b[3],cfgb_mirn_b[2],cfgb_mirn_b[1]
*.ipin cfgb_mirp_b[6],cfgb_mirp_b[5],cfgb_mirp_b[4],cfgb_mirp_b[3],cfgb_mirp_b[2],cfgb_mirp_b[1]
*.ipin cfgb_dpn_inm[3],cfgb_dpn_inm[2],cfgb_dpn_inm[1]
*.ipin
*+ cfgb_dpn_outm[6],cfgb_dpn_outm[5],cfgb_dpn_outm[4],cfgb_dpn_outm[3],cfgb_dpn_outm[2],cfgb_dpn_outm[1]
*.ipin cfgb_dpp_inm[3],cfgb_dpp_inm[2],cfgb_dpp_inm[1]
*.ipin
*+ cfgb_dpp_outm[6],cfgb_dpp_outm[5],cfgb_dpp_outm[4],cfgb_dpp_outm[3],cfgb_dpp_outm[2],cfgb_dpp_outm[1]
*.ipin
*+ cfgb_nfetb_d[6],cfgb_nfetb_d[5],cfgb_nfetb_d[4],cfgb_nfetb_d[3],cfgb_nfetb_d[2],cfgb_nfetb_d[1]
*.ipin
*+ cfgb_nfetb_g[6],cfgb_nfetb_g[5],cfgb_nfetb_g[4],cfgb_nfetb_g[3],cfgb_nfetb_g[2],cfgb_nfetb_g[1]
*.ipin
*+ cfgb_nfetb_s[6],cfgb_nfetb_s[5],cfgb_nfetb_s[4],cfgb_nfetb_s[3],cfgb_nfetb_s[2],cfgb_nfetb_s[1]
*.ipin
*+ cfgb_pfetb_d[6],cfgb_pfetb_d[5],cfgb_pfetb_d[4],cfgb_pfetb_d[3],cfgb_pfetb_d[2],cfgb_pfetb_d[1]
*.ipin
*+ cfgb_pfetb_g[6],cfgb_pfetb_g[5],cfgb_pfetb_g[4],cfgb_pfetb_g[3],cfgb_pfetb_g[2],cfgb_pfetb_g[1]
*.ipin
*+ cfgb_pfetb_s[6],cfgb_pfetb_s[5],cfgb_pfetb_s[4],cfgb_pfetb_s[3],cfgb_pfetb_s[2],cfgb_pfetb_s[1]
*.ipin ibias
*.ipin
*+ cfg_bus_short[6],cfg_bus_short[5],cfg_bus_short[4],cfg_bus_short[3],cfg_bus_short[2],cfg_bus_short[1]
*.ipin ctrl_otan_tail[1],ctrl_otan_tail[0]
*.ipin ctrl_otan_diode
*.ipin ctrl_mirn_a[1],ctrl_mirn_a[0]
*.ipin ctrl_mirn_b[1],ctrl_mirn_b[0]
*.ipin ctrl_mirp_a[1],ctrl_mirp_a[0]
*.ipin ctrl_mirp_b[1],ctrl_mirp_b[0]
*.ipin ctrl_dpn_tail[1],ctrl_dpn_tail[0]
*.ipin ctrl_dpn_source
*.ipin ctrl_dpp_tail[1],ctrl_dpp_tail[0]
*.ipin ctrl_dpp_source
*.ipin ctrl_nfeta_width[1],ctrl_nfeta_width[0]
*.ipin ctrl_nfeta_source
*.ipin ctrl_nfetb_width[1],ctrl_nfetb_width[0]
*.ipin ctrl_nfetb_source
*.ipin ctrl_pfeta_width[1],ctrl_pfeta_width[0]
*.ipin ctrl_pfeta_source
*.ipin ctrl_pfetb_width[1],ctrl_pfetb_width[0]
*.ipin ctrl_pfetb_source
*.iopin VAPWR
*.iopin VDPWR
*.iopin VGND
*.iopin bus_A[5],bus_A[4],bus_A[3],bus_A[2],bus_A[1]
*.ipin cfg_bus_ext[5],cfg_bus_ext[4],cfg_bus_ext[3],cfg_bus_ext[2],cfg_bus_ext[1]
x2 VAPWR VDPWR ibias ibias_p xpt_mirn_a xpt_mirn_b ctrl_mirn_a[1] ctrl_mirn_a[0] ctrl_mirn_b[1]
+ ctrl_mirn_b[0] VGND mirror_n
x10[6] VGND VDPWR VAPWR cfga_vapwr[6] VAPWR bus_A_int[6] tt_asw_3v3
x10[5] VGND VDPWR VAPWR cfga_vapwr[5] VAPWR bus_A_int[5] tt_asw_3v3
x10[4] VGND VDPWR VAPWR cfga_vapwr[4] VAPWR bus_A_int[4] tt_asw_3v3
x10[3] VGND VDPWR VAPWR cfga_vapwr[3] VAPWR bus_A_int[3] tt_asw_3v3
x10[2] VGND VDPWR VAPWR cfga_vapwr[2] VAPWR bus_A_int[2] tt_asw_3v3
x10[1] VGND VDPWR VAPWR cfga_vapwr[1] VAPWR bus_A_int[1] tt_asw_3v3
x11[6] VGND VDPWR VAPWR cfga_vgnd[6] VGND bus_A_int[6] tt_asw_3v3
x11[5] VGND VDPWR VAPWR cfga_vgnd[5] VGND bus_A_int[5] tt_asw_3v3
x11[4] VGND VDPWR VAPWR cfga_vgnd[4] VGND bus_A_int[4] tt_asw_3v3
x11[3] VGND VDPWR VAPWR cfga_vgnd[3] VGND bus_A_int[3] tt_asw_3v3
x11[2] VGND VDPWR VAPWR cfga_vgnd[2] VGND bus_A_int[2] tt_asw_3v3
x11[1] VGND VDPWR VAPWR cfga_vgnd[1] VGND bus_A_int[1] tt_asw_3v3
x12[3] VGND VDPWR VAPWR cfga_otan_inp[3] xpt_otan_inp bus_A_int[3] tt_asw_3v3
x12[2] VGND VDPWR VAPWR cfga_otan_inp[2] xpt_otan_inp bus_A_int[2] tt_asw_3v3
x12[1] VGND VDPWR VAPWR cfga_otan_inp[1] xpt_otan_inp bus_A_int[1] tt_asw_3v3
x13[6] VGND VDPWR VAPWR cfga_otan_out[6] xpt_otan_out bus_A_int[6] tt_asw_3v3
x13[5] VGND VDPWR VAPWR cfga_otan_out[5] xpt_otan_out bus_A_int[5] tt_asw_3v3
x13[4] VGND VDPWR VAPWR cfga_otan_out[4] xpt_otan_out bus_A_int[4] tt_asw_3v3
x13[3] VGND VDPWR VAPWR cfga_otan_out[3] xpt_otan_out bus_A_int[3] tt_asw_3v3
x13[2] VGND VDPWR VAPWR cfga_otan_out[2] xpt_otan_out bus_A_int[2] tt_asw_3v3
x13[1] VGND VDPWR VAPWR cfga_otan_out[1] xpt_otan_out bus_A_int[1] tt_asw_3v3
x14[6] VGND VDPWR VAPWR cfga_mirn_a[6] xpt_mirn_a bus_A_int[6] tt_asw_3v3
x14[5] VGND VDPWR VAPWR cfga_mirn_a[5] xpt_mirn_a bus_A_int[5] tt_asw_3v3
x14[4] VGND VDPWR VAPWR cfga_mirn_a[4] xpt_mirn_a bus_A_int[4] tt_asw_3v3
x14[3] VGND VDPWR VAPWR cfga_mirn_a[3] xpt_mirn_a bus_A_int[3] tt_asw_3v3
x14[2] VGND VDPWR VAPWR cfga_mirn_a[2] xpt_mirn_a bus_A_int[2] tt_asw_3v3
x14[1] VGND VDPWR VAPWR cfga_mirn_a[1] xpt_mirn_a bus_A_int[1] tt_asw_3v3
x15[6] VGND VDPWR VAPWR cfga_mirp_a[6] xpt_mirp_a bus_A_int[6] tt_asw_3v3
x15[5] VGND VDPWR VAPWR cfga_mirp_a[5] xpt_mirp_a bus_A_int[5] tt_asw_3v3
x15[4] VGND VDPWR VAPWR cfga_mirp_a[4] xpt_mirp_a bus_A_int[4] tt_asw_3v3
x15[3] VGND VDPWR VAPWR cfga_mirp_a[3] xpt_mirp_a bus_A_int[3] tt_asw_3v3
x15[2] VGND VDPWR VAPWR cfga_mirp_a[2] xpt_mirp_a bus_A_int[2] tt_asw_3v3
x15[1] VGND VDPWR VAPWR cfga_mirp_a[1] xpt_mirp_a bus_A_int[1] tt_asw_3v3
x16[3] VGND VDPWR VAPWR cfga_dpn_inp[3] xpt_dpn_inp bus_A_int[3] tt_asw_3v3
x16[2] VGND VDPWR VAPWR cfga_dpn_inp[2] xpt_dpn_inp bus_A_int[2] tt_asw_3v3
x16[1] VGND VDPWR VAPWR cfga_dpn_inp[1] xpt_dpn_inp bus_A_int[1] tt_asw_3v3
x17[6] VGND VDPWR VAPWR cfga_dpn_outp[6] xpt_dpn_outp bus_A_int[6] tt_asw_3v3
x17[5] VGND VDPWR VAPWR cfga_dpn_outp[5] xpt_dpn_outp bus_A_int[5] tt_asw_3v3
x17[4] VGND VDPWR VAPWR cfga_dpn_outp[4] xpt_dpn_outp bus_A_int[4] tt_asw_3v3
x17[3] VGND VDPWR VAPWR cfga_dpn_outp[3] xpt_dpn_outp bus_A_int[3] tt_asw_3v3
x17[2] VGND VDPWR VAPWR cfga_dpn_outp[2] xpt_dpn_outp bus_A_int[2] tt_asw_3v3
x17[1] VGND VDPWR VAPWR cfga_dpn_outp[1] xpt_dpn_outp bus_A_int[1] tt_asw_3v3
x18[3] VGND VDPWR VAPWR cfga_dpp_inp[3] xpt_dpp_inp bus_A_int[3] tt_asw_3v3
x18[2] VGND VDPWR VAPWR cfga_dpp_inp[2] xpt_dpp_inp bus_A_int[2] tt_asw_3v3
x18[1] VGND VDPWR VAPWR cfga_dpp_inp[1] xpt_dpp_inp bus_A_int[1] tt_asw_3v3
x19[6] VGND VDPWR VAPWR cfga_dpp_outp[6] xpt_dpp_outp bus_A_int[6] tt_asw_3v3
x19[5] VGND VDPWR VAPWR cfga_dpp_outp[5] xpt_dpp_outp bus_A_int[5] tt_asw_3v3
x19[4] VGND VDPWR VAPWR cfga_dpp_outp[4] xpt_dpp_outp bus_A_int[4] tt_asw_3v3
x19[3] VGND VDPWR VAPWR cfga_dpp_outp[3] xpt_dpp_outp bus_A_int[3] tt_asw_3v3
x19[2] VGND VDPWR VAPWR cfga_dpp_outp[2] xpt_dpp_outp bus_A_int[2] tt_asw_3v3
x19[1] VGND VDPWR VAPWR cfga_dpp_outp[1] xpt_dpp_outp bus_A_int[1] tt_asw_3v3
x20[6] VGND VDPWR VAPWR cfga_nfeta_d[6] xpt_nfeta_d bus_A_int[6] tt_asw_3v3
x20[5] VGND VDPWR VAPWR cfga_nfeta_d[5] xpt_nfeta_d bus_A_int[5] tt_asw_3v3
x20[4] VGND VDPWR VAPWR cfga_nfeta_d[4] xpt_nfeta_d bus_A_int[4] tt_asw_3v3
x20[3] VGND VDPWR VAPWR cfga_nfeta_d[3] xpt_nfeta_d bus_A_int[3] tt_asw_3v3
x20[2] VGND VDPWR VAPWR cfga_nfeta_d[2] xpt_nfeta_d bus_A_int[2] tt_asw_3v3
x20[1] VGND VDPWR VAPWR cfga_nfeta_d[1] xpt_nfeta_d bus_A_int[1] tt_asw_3v3
x21[6] VGND VDPWR VAPWR cfga_nfeta_g[6] xpt_nfeta_g bus_A_int[6] tt_asw_3v3
x21[5] VGND VDPWR VAPWR cfga_nfeta_g[5] xpt_nfeta_g bus_A_int[5] tt_asw_3v3
x21[4] VGND VDPWR VAPWR cfga_nfeta_g[4] xpt_nfeta_g bus_A_int[4] tt_asw_3v3
x21[3] VGND VDPWR VAPWR cfga_nfeta_g[3] xpt_nfeta_g bus_A_int[3] tt_asw_3v3
x21[2] VGND VDPWR VAPWR cfga_nfeta_g[2] xpt_nfeta_g bus_A_int[2] tt_asw_3v3
x21[1] VGND VDPWR VAPWR cfga_nfeta_g[1] xpt_nfeta_g bus_A_int[1] tt_asw_3v3
x22[6] VGND VDPWR VAPWR cfga_nfeta_s[6] xpt_nfeta_s bus_A_int[6] tt_asw_3v3
x22[5] VGND VDPWR VAPWR cfga_nfeta_s[5] xpt_nfeta_s bus_A_int[5] tt_asw_3v3
x22[4] VGND VDPWR VAPWR cfga_nfeta_s[4] xpt_nfeta_s bus_A_int[4] tt_asw_3v3
x22[3] VGND VDPWR VAPWR cfga_nfeta_s[3] xpt_nfeta_s bus_A_int[3] tt_asw_3v3
x22[2] VGND VDPWR VAPWR cfga_nfeta_s[2] xpt_nfeta_s bus_A_int[2] tt_asw_3v3
x22[1] VGND VDPWR VAPWR cfga_nfeta_s[1] xpt_nfeta_s bus_A_int[1] tt_asw_3v3
x23[6] VGND VDPWR VAPWR cfga_pfeta_d[6] xpt_pfeta_d bus_A_int[6] tt_asw_3v3
x23[5] VGND VDPWR VAPWR cfga_pfeta_d[5] xpt_pfeta_d bus_A_int[5] tt_asw_3v3
x23[4] VGND VDPWR VAPWR cfga_pfeta_d[4] xpt_pfeta_d bus_A_int[4] tt_asw_3v3
x23[3] VGND VDPWR VAPWR cfga_pfeta_d[3] xpt_pfeta_d bus_A_int[3] tt_asw_3v3
x23[2] VGND VDPWR VAPWR cfga_pfeta_d[2] xpt_pfeta_d bus_A_int[2] tt_asw_3v3
x23[1] VGND VDPWR VAPWR cfga_pfeta_d[1] xpt_pfeta_d bus_A_int[1] tt_asw_3v3
x24[6] VGND VDPWR VAPWR cfga_pfeta_g[6] xpt_pfeta_g bus_A_int[6] tt_asw_3v3
x24[5] VGND VDPWR VAPWR cfga_pfeta_g[5] xpt_pfeta_g bus_A_int[5] tt_asw_3v3
x24[4] VGND VDPWR VAPWR cfga_pfeta_g[4] xpt_pfeta_g bus_A_int[4] tt_asw_3v3
x24[3] VGND VDPWR VAPWR cfga_pfeta_g[3] xpt_pfeta_g bus_A_int[3] tt_asw_3v3
x24[2] VGND VDPWR VAPWR cfga_pfeta_g[2] xpt_pfeta_g bus_A_int[2] tt_asw_3v3
x24[1] VGND VDPWR VAPWR cfga_pfeta_g[1] xpt_pfeta_g bus_A_int[1] tt_asw_3v3
x25[6] VGND VDPWR VAPWR cfga_pfeta_s[6] xpt_pfeta_s bus_A_int[6] tt_asw_3v3
x25[5] VGND VDPWR VAPWR cfga_pfeta_s[5] xpt_pfeta_s bus_A_int[5] tt_asw_3v3
x25[4] VGND VDPWR VAPWR cfga_pfeta_s[4] xpt_pfeta_s bus_A_int[4] tt_asw_3v3
x25[3] VGND VDPWR VAPWR cfga_pfeta_s[3] xpt_pfeta_s bus_A_int[3] tt_asw_3v3
x25[2] VGND VDPWR VAPWR cfga_pfeta_s[2] xpt_pfeta_s bus_A_int[2] tt_asw_3v3
x25[1] VGND VDPWR VAPWR cfga_pfeta_s[1] xpt_pfeta_s bus_A_int[1] tt_asw_3v3
x28[3] VGND VDPWR VAPWR cfgb_otan_inm[3] xpt_otan_inm bus_B_int[3] tt_asw_3v3
x28[2] VGND VDPWR VAPWR cfgb_otan_inm[2] xpt_otan_inm bus_B_int[2] tt_asw_3v3
x28[1] VGND VDPWR VAPWR cfgb_otan_inm[1] xpt_otan_inm bus_B_int[1] tt_asw_3v3
x30[6] VGND VDPWR VAPWR cfgb_mirn_b[6] xpt_mirn_b bus_B_int[6] tt_asw_3v3
x30[5] VGND VDPWR VAPWR cfgb_mirn_b[5] xpt_mirn_b bus_B_int[5] tt_asw_3v3
x30[4] VGND VDPWR VAPWR cfgb_mirn_b[4] xpt_mirn_b bus_B_int[4] tt_asw_3v3
x30[3] VGND VDPWR VAPWR cfgb_mirn_b[3] xpt_mirn_b bus_B_int[3] tt_asw_3v3
x30[2] VGND VDPWR VAPWR cfgb_mirn_b[2] xpt_mirn_b bus_B_int[2] tt_asw_3v3
x30[1] VGND VDPWR VAPWR cfgb_mirn_b[1] xpt_mirn_b bus_B_int[1] tt_asw_3v3
x31[6] VGND VDPWR VAPWR cfgb_mirp_b[6] xpt_mirp_b bus_B_int[6] tt_asw_3v3
x31[5] VGND VDPWR VAPWR cfgb_mirp_b[5] xpt_mirp_b bus_B_int[5] tt_asw_3v3
x31[4] VGND VDPWR VAPWR cfgb_mirp_b[4] xpt_mirp_b bus_B_int[4] tt_asw_3v3
x31[3] VGND VDPWR VAPWR cfgb_mirp_b[3] xpt_mirp_b bus_B_int[3] tt_asw_3v3
x31[2] VGND VDPWR VAPWR cfgb_mirp_b[2] xpt_mirp_b bus_B_int[2] tt_asw_3v3
x31[1] VGND VDPWR VAPWR cfgb_mirp_b[1] xpt_mirp_b bus_B_int[1] tt_asw_3v3
x32[3] VGND VDPWR VAPWR cfgb_dpn_inm[3] xpt_dpn_inm bus_B_int[3] tt_asw_3v3
x32[2] VGND VDPWR VAPWR cfgb_dpn_inm[2] xpt_dpn_inm bus_B_int[2] tt_asw_3v3
x32[1] VGND VDPWR VAPWR cfgb_dpn_inm[1] xpt_dpn_inm bus_B_int[1] tt_asw_3v3
x33[6] VGND VDPWR VAPWR cfgb_dpn_outm[6] xpt_dpn_outm bus_B_int[6] tt_asw_3v3
x33[5] VGND VDPWR VAPWR cfgb_dpn_outm[5] xpt_dpn_outm bus_B_int[5] tt_asw_3v3
x33[4] VGND VDPWR VAPWR cfgb_dpn_outm[4] xpt_dpn_outm bus_B_int[4] tt_asw_3v3
x33[3] VGND VDPWR VAPWR cfgb_dpn_outm[3] xpt_dpn_outm bus_B_int[3] tt_asw_3v3
x33[2] VGND VDPWR VAPWR cfgb_dpn_outm[2] xpt_dpn_outm bus_B_int[2] tt_asw_3v3
x33[1] VGND VDPWR VAPWR cfgb_dpn_outm[1] xpt_dpn_outm bus_B_int[1] tt_asw_3v3
x34[3] VGND VDPWR VAPWR cfgb_dpp_inm[3] xpt_dpp_inm bus_B_int[3] tt_asw_3v3
x34[2] VGND VDPWR VAPWR cfgb_dpp_inm[2] xpt_dpp_inm bus_B_int[2] tt_asw_3v3
x34[1] VGND VDPWR VAPWR cfgb_dpp_inm[1] xpt_dpp_inm bus_B_int[1] tt_asw_3v3
x35[6] VGND VDPWR VAPWR cfgb_dpp_outm[6] xpt_dpp_outm bus_B_int[6] tt_asw_3v3
x35[5] VGND VDPWR VAPWR cfgb_dpp_outm[5] xpt_dpp_outm bus_B_int[5] tt_asw_3v3
x35[4] VGND VDPWR VAPWR cfgb_dpp_outm[4] xpt_dpp_outm bus_B_int[4] tt_asw_3v3
x35[3] VGND VDPWR VAPWR cfgb_dpp_outm[3] xpt_dpp_outm bus_B_int[3] tt_asw_3v3
x35[2] VGND VDPWR VAPWR cfgb_dpp_outm[2] xpt_dpp_outm bus_B_int[2] tt_asw_3v3
x35[1] VGND VDPWR VAPWR cfgb_dpp_outm[1] xpt_dpp_outm bus_B_int[1] tt_asw_3v3
x36[6] VGND VDPWR VAPWR cfgb_nfetb_d[6] xpt_nfetb_d bus_B_int[6] tt_asw_3v3
x36[5] VGND VDPWR VAPWR cfgb_nfetb_d[5] xpt_nfetb_d bus_B_int[5] tt_asw_3v3
x36[4] VGND VDPWR VAPWR cfgb_nfetb_d[4] xpt_nfetb_d bus_B_int[4] tt_asw_3v3
x36[3] VGND VDPWR VAPWR cfgb_nfetb_d[3] xpt_nfetb_d bus_B_int[3] tt_asw_3v3
x36[2] VGND VDPWR VAPWR cfgb_nfetb_d[2] xpt_nfetb_d bus_B_int[2] tt_asw_3v3
x36[1] VGND VDPWR VAPWR cfgb_nfetb_d[1] xpt_nfetb_d bus_B_int[1] tt_asw_3v3
x37[6] VGND VDPWR VAPWR cfgb_nfetb_g[6] xpt_nfetb_g bus_B_int[6] tt_asw_3v3
x37[5] VGND VDPWR VAPWR cfgb_nfetb_g[5] xpt_nfetb_g bus_B_int[5] tt_asw_3v3
x37[4] VGND VDPWR VAPWR cfgb_nfetb_g[4] xpt_nfetb_g bus_B_int[4] tt_asw_3v3
x37[3] VGND VDPWR VAPWR cfgb_nfetb_g[3] xpt_nfetb_g bus_B_int[3] tt_asw_3v3
x37[2] VGND VDPWR VAPWR cfgb_nfetb_g[2] xpt_nfetb_g bus_B_int[2] tt_asw_3v3
x37[1] VGND VDPWR VAPWR cfgb_nfetb_g[1] xpt_nfetb_g bus_B_int[1] tt_asw_3v3
x38[6] VGND VDPWR VAPWR cfgb_nfetb_s[6] xpt_nfetb_s bus_B_int[6] tt_asw_3v3
x38[5] VGND VDPWR VAPWR cfgb_nfetb_s[5] xpt_nfetb_s bus_B_int[5] tt_asw_3v3
x38[4] VGND VDPWR VAPWR cfgb_nfetb_s[4] xpt_nfetb_s bus_B_int[4] tt_asw_3v3
x38[3] VGND VDPWR VAPWR cfgb_nfetb_s[3] xpt_nfetb_s bus_B_int[3] tt_asw_3v3
x38[2] VGND VDPWR VAPWR cfgb_nfetb_s[2] xpt_nfetb_s bus_B_int[2] tt_asw_3v3
x38[1] VGND VDPWR VAPWR cfgb_nfetb_s[1] xpt_nfetb_s bus_B_int[1] tt_asw_3v3
x39[6] VGND VDPWR VAPWR cfgb_pfetb_d[6] xpt_pfetb_d bus_B_int[6] tt_asw_3v3
x39[5] VGND VDPWR VAPWR cfgb_pfetb_d[5] xpt_pfetb_d bus_B_int[5] tt_asw_3v3
x39[4] VGND VDPWR VAPWR cfgb_pfetb_d[4] xpt_pfetb_d bus_B_int[4] tt_asw_3v3
x39[3] VGND VDPWR VAPWR cfgb_pfetb_d[3] xpt_pfetb_d bus_B_int[3] tt_asw_3v3
x39[2] VGND VDPWR VAPWR cfgb_pfetb_d[2] xpt_pfetb_d bus_B_int[2] tt_asw_3v3
x39[1] VGND VDPWR VAPWR cfgb_pfetb_d[1] xpt_pfetb_d bus_B_int[1] tt_asw_3v3
x40[6] VGND VDPWR VAPWR cfgb_pfetb_g[6] xpt_pfetb_g bus_B_int[6] tt_asw_3v3
x40[5] VGND VDPWR VAPWR cfgb_pfetb_g[5] xpt_pfetb_g bus_B_int[5] tt_asw_3v3
x40[4] VGND VDPWR VAPWR cfgb_pfetb_g[4] xpt_pfetb_g bus_B_int[4] tt_asw_3v3
x40[3] VGND VDPWR VAPWR cfgb_pfetb_g[3] xpt_pfetb_g bus_B_int[3] tt_asw_3v3
x40[2] VGND VDPWR VAPWR cfgb_pfetb_g[2] xpt_pfetb_g bus_B_int[2] tt_asw_3v3
x40[1] VGND VDPWR VAPWR cfgb_pfetb_g[1] xpt_pfetb_g bus_B_int[1] tt_asw_3v3
x41[6] VGND VDPWR VAPWR cfgb_pfetb_s[6] xpt_pfetb_s bus_B_int[6] tt_asw_3v3
x41[5] VGND VDPWR VAPWR cfgb_pfetb_s[5] xpt_pfetb_s bus_B_int[5] tt_asw_3v3
x41[4] VGND VDPWR VAPWR cfgb_pfetb_s[4] xpt_pfetb_s bus_B_int[4] tt_asw_3v3
x41[3] VGND VDPWR VAPWR cfgb_pfetb_s[3] xpt_pfetb_s bus_B_int[3] tt_asw_3v3
x41[2] VGND VDPWR VAPWR cfgb_pfetb_s[2] xpt_pfetb_s bus_B_int[2] tt_asw_3v3
x41[1] VGND VDPWR VAPWR cfgb_pfetb_s[1] xpt_pfetb_s bus_B_int[1] tt_asw_3v3
x42[6] VGND VDPWR VAPWR cfg_bus_short[6] bus_A_int[6] bus_B_int[6] tt_asw_3v3
x42[5] VGND VDPWR VAPWR cfg_bus_short[5] bus_A_int[5] bus_B_int[5] tt_asw_3v3
x42[4] VGND VDPWR VAPWR cfg_bus_short[4] bus_A_int[4] bus_B_int[4] tt_asw_3v3
x42[3] VGND VDPWR VAPWR cfg_bus_short[3] bus_A_int[3] bus_B_int[3] tt_asw_3v3
x42[2] VGND VDPWR VAPWR cfg_bus_short[2] bus_A_int[2] bus_B_int[2] tt_asw_3v3
x42[1] VGND VDPWR VAPWR cfg_bus_short[1] bus_A_int[1] bus_B_int[1] tt_asw_3v3
x1 VAPWR VDPWR xpt_otan_inp xpt_otan_out xpt_otan_inm ctrl_otan_tail[1] ctrl_otan_tail[0]
+ ctrl_otan_diode ibias VGND ota_n
x3 VAPWR VDPWR ibias_p xpt_mirp_a xpt_mirp_b ctrl_mirp_a[1] ctrl_mirp_a[0] ctrl_mirp_b[1]
+ ctrl_mirp_b[0] VGND mirror_p
x4 VAPWR VDPWR xpt_dpn_outp xpt_dpn_outm xpt_dpn_inp xpt_dpn_inm ctrl_dpn_tail[1] ctrl_dpn_tail[0]
+ ctrl_dpn_source ibias VGND diff_n
x5 VAPWR VDPWR xpt_dpp_outp xpt_dpp_outm xpt_dpp_inp xpt_dpp_inm ctrl_dpp_tail[1] ctrl_dpp_tail[0]
+ ctrl_dpp_source ibias_p VGND diff_p
x6 VAPWR VDPWR xpt_nfeta_d xpt_nfeta_g xpt_nfeta_s ctrl_nfeta_source ctrl_nfeta_width[1]
+ ctrl_nfeta_width[0] VGND nmos_prog
x7 VAPWR VDPWR xpt_nfetb_d xpt_nfetb_g xpt_nfetb_s ctrl_nfetb_source ctrl_nfetb_width[1]
+ ctrl_nfetb_width[0] VGND nmos_prog
x8 VAPWR VDPWR xpt_pfeta_s xpt_pfeta_g xpt_pfeta_d ctrl_pfeta_source ctrl_pfeta_width[1]
+ ctrl_pfeta_width[0] VGND pmos_prog
x9 VAPWR VDPWR xpt_pfetb_s xpt_pfetb_g xpt_pfetb_d ctrl_pfetb_source ctrl_pfetb_width[1]
+ ctrl_pfetb_width[0] VGND pmos_prog
x1[5] VGND VDPWR VAPWR cfg_bus_ext[5] bus_A[5] bus_A_int[5] tt_asw_3v3
x1[4] VGND VDPWR VAPWR cfg_bus_ext[4] bus_A[4] bus_A_int[4] tt_asw_3v3
x1[3] VGND VDPWR VAPWR cfg_bus_ext[3] bus_A[3] bus_A_int[3] tt_asw_3v3
x1[2] VGND VDPWR VAPWR cfg_bus_ext[2] bus_A[2] bus_A_int[2] tt_asw_3v3
x1[1] VGND VDPWR VAPWR cfg_bus_ext[1] bus_A[1] bus_A_int[1] tt_asw_3v3
.ends


* expanding   symbol:  mirror_n.sym # of pins=9
** sym_path: /foss/designs/ttsky25a_minimosbius/xschem/mirror_n.sym
** sch_path: /foss/designs/ttsky25a_minimosbius/xschem/mirror_n.sch
.subckt mirror_n VAPWR VDPWR ibias iout_fixed iout_1 iout_2 ictrl_1[1] ictrl_1[0] ictrl_2[1]
+ ictrl_2[0] GND
*.iopin ibias
*.iopin iout_fixed
*.iopin iout_1
*.ipin ictrl_1[1],ictrl_1[0]
*.ipin ictrl_2[1],ictrl_2[0]
*.iopin iout_2
*.iopin VAPWR
*.iopin VDPWR
*.iopin GND
XM1 ibias ibias GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=10 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 iout_fixed ibias GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=10 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 i1_1x ibias GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=10 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 iout_1 ibias GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=10 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 i1_2x ibias GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=20 nf=4 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x4 GND VDPWR VAPWR ictrl_1[0] i1_1x iout_1 tt_asw_3v3
x5 GND VDPWR VAPWR ictrl_1[1] i1_2x iout_1 tt_asw_3v3
XM14 i2_1x ibias GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=10 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM16 iout_2 ibias GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=10 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18 i2_2x ibias GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=20 nf=4 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x1 GND VDPWR VAPWR ictrl_2[0] i2_1x iout_2 tt_asw_3v3
x2 GND VDPWR VAPWR ictrl_2[1] i2_2x iout_2 tt_asw_3v3
XM4 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=20 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  pad_model.sym # of pins=3
** sym_path: /foss/designs/ttsky25a_minimosbius/xschem/pad_model.sym
** sch_path: /foss/designs/ttsky25a_minimosbius/xschem/pad_model.sch
.subckt pad_model VGND pin mod
*.iopin pin
*.iopin mod
*.iopin VGND
XM1 net3 VAPWR mod VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=60 nf=12 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net3 VGND mod VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=180 nf=18 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
C1 pin VGND 2p m=1
V1 VAPWR VGND 3.3
.save i(v1)
R1 net1 pin 1 m=1
L1 net2 net1 1n m=1
C2 net2 VGND 3p m=1
R2 net3 net2 50 m=1
C3 mod VGND 250f m=1
XM3 net3 VGND VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=60 nf=12 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=15 m=15
XM4 net3 VAPWR VGND VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=180 nf=18 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=15 m=15
.ends


* expanding   symbol:  diff_n.sym # of pins=10
** sym_path: /foss/designs/ttsky25a_minimosbius/xschem/diff_n.sym
** sch_path: /foss/designs/ttsky25a_minimosbius/xschem/diff_n.sch
.subckt diff_n VAPWR VDPWR outp outm inp inm ctrl_tail[1] ctrl_tail[0] ctrl_source vbias GND
*.iopin vbias
*.ipin ctrl_tail[1],ctrl_tail[0]
*.iopin VAPWR
*.iopin VDPWR
*.iopin GND
*.ipin ctrl_source
*.ipin inp
*.ipin inm
*.iopin outp
*.iopin outm
XM1 outp inp itail itail sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=40 nf=8 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 outm inm itail itail sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=40 nf=8 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 itail_1x vbias GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=20 nf=4 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 itail vbias GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=20 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 itail_2x vbias GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=40 nf=8 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x4 GND VDPWR VAPWR ctrl_tail[0] itail_1x itail tt_asw_3v3
x5 GND VDPWR VAPWR ctrl_tail[1] itail_2x itail tt_asw_3v3
x1 GND VDPWR VAPWR ctrl_source itail GND tt_asw_3v3
XM3 itail itail itail itail sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  tt_asw_3v3.sym # of pins=6
** sym_path: /foss/designs/ttsky25a_minimosbius/xschem/tt_asw_3v3.sym
** sch_path: /foss/designs/ttsky25a_minimosbius/xschem/tt_asw_3v3.sch
.subckt tt_asw_3v3 VGND VDPWR VAPWR ctrl mod bus
*.iopin mod
*.iopin bus
*.ipin ctrl
*.iopin VGND
*.iopin VDPWR
*.iopin VAPWR
XM1 tgon_n net2 VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 tgon_n net2 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 tgon net1 VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 tgon net1 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 bus tgon_n mod VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=180 nf=18 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 bus tgon mod VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=60 nf=12 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 ctrl_n ctrl VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 ctrl_n ctrl VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net1 ctrl VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 net2 ctrl_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 net1 net2 net3 VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 net2 net1 net4 VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 net3 net1 VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 net4 net2 VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  ota_n.sym # of pins=9
** sym_path: /foss/designs/ttsky25a_minimosbius/xschem/ota_n.sym
** sch_path: /foss/designs/ttsky25a_minimosbius/xschem/ota_n.sch
.subckt ota_n VAPWR VDPWR inp out inm ctrl_tail[1] ctrl_tail[0] ctrl_diode vbias GND
*.iopin vbias
*.ipin ctrl_tail[1],ctrl_tail[0]
*.iopin VAPWR
*.iopin VDPWR
*.iopin GND
*.ipin ctrl_diode
*.ipin inp
*.ipin inm
*.opin out
XM1 outb outb VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=1 W=60 nf=12 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 out out_gate VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=1 W=60 nf=12 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x2 GND VDPWR VAPWR ctrl_diode_b outb out_gate tt_asw_3v3
x3 GND VDPWR VAPWR ctrl_diode out out_gate tt_asw_3v3
XM7 ctrl_diode_b ctrl_diode GND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 ctrl_diode_b ctrl_diode VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 VAPWR VAPWR VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=1 W=10 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 outb inp itail itail sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=40 nf=8 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 out inm itail itail sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=40 nf=8 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 itail_1x vbias GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=20 nf=4 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 itail vbias GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=20 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 itail_2x vbias GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=40 nf=8 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x4 GND VDPWR VAPWR ctrl_tail[0] itail_1x itail tt_asw_3v3
x5 GND VDPWR VAPWR ctrl_tail[1] itail_2x itail tt_asw_3v3
.ends


* expanding   symbol:  mirror_p.sym # of pins=8
** sym_path: /foss/designs/ttsky25a_minimosbius/xschem/mirror_p.sym
** sch_path: /foss/designs/ttsky25a_minimosbius/xschem/mirror_p.sch
.subckt mirror_p VAPWR VDPWR ibias iout_1 iout_2 ictrl_1[1] ictrl_1[0] ictrl_2[1] ictrl_2[0] GND
*.iopin ibias
*.iopin iout_1
*.ipin ictrl_1[1],ictrl_1[0]
*.ipin ictrl_2[1],ictrl_2[0]
*.iopin iout_2
*.iopin VAPWR
*.iopin VDPWR
*.iopin GND
x4 GND VDPWR VAPWR ictrl_1[0] i1_1x iout_1 tt_asw_3v3
x5 GND VDPWR VAPWR ictrl_1[1] i1_2x iout_1 tt_asw_3v3
x1 GND VDPWR VAPWR ictrl_2[0] i2_1x iout_2 tt_asw_3v3
x2 GND VDPWR VAPWR ictrl_2[1] i2_2x iout_2 tt_asw_3v3
XM3 iout_1 ibias VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=1 W=30 nf=6 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 ibias ibias VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=1 W=30 nf=6 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 i1_1x ibias VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=1 W=30 nf=6 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 i1_2x ibias VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=1 W=60 nf=12 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 iout_2 ibias VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=1 W=30 nf=6 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 i2_1x ibias VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=1 W=30 nf=6 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 i2_2x ibias VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=1 W=60 nf=12 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  diff_p.sym # of pins=10
** sym_path: /foss/designs/ttsky25a_minimosbius/xschem/diff_p.sym
** sch_path: /foss/designs/ttsky25a_minimosbius/xschem/diff_p.sch
.subckt diff_p VAPWR VDPWR outp outm inp inm ctrl_tail[1] ctrl_tail[0] ctrl_source vbias GND
*.iopin vbias
*.ipin ctrl_tail[1],ctrl_tail[0]
*.iopin VAPWR
*.iopin VDPWR
*.iopin GND
*.ipin ctrl_source
*.ipin inp
*.ipin inm
*.iopin outp
*.iopin outm
x4 GND VDPWR VAPWR ctrl_tail[0] itail_1x itail tt_asw_3v3
x5 GND VDPWR VAPWR ctrl_tail[1] itail_2x itail tt_asw_3v3
x1 GND VDPWR VAPWR ctrl_source itail VAPWR tt_asw_3v3
XM3 outp inp itail itail sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=120 nf=24 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 outm inm itail itail sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=120 nf=24 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 itail vbias VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=1 W=60 nf=12 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 itail_1x vbias VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=1 W=60 nf=12 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 itail_2x vbias VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=1 W=120 nf=24 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  nmos_prog.sym # of pins=8
** sym_path: /foss/designs/ttsky25a_minimosbius/xschem/nmos_prog.sym
** sch_path: /foss/designs/ttsky25a_minimosbius/xschem/nmos_prog.sch
.subckt nmos_prog VAPWR VDPWR Vd Vg Vs ctrl_source ctrl_width[1] ctrl_width[0] GND
*.ipin ctrl_width[1],ctrl_width[0]
*.iopin Vs
*.iopin Vg
*.iopin Vd
*.iopin VAPWR
*.iopin VDPWR
*.iopin GND
*.ipin ctrl_source
XM1 Vd Vg Vs Vs sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vd_1x Vg Vs Vs sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vd_2x Vg Vs Vs sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
x1 GND VDPWR VAPWR ctrl_width[0] Vd_1x Vd tt_asw_3v3
x2 GND VDPWR VAPWR ctrl_width[1] Vd_2x Vd tt_asw_3v3
x3 GND VDPWR VAPWR ctrl_source Vs GND tt_asw_3v3
XM4 Vs Vs Vs Vs sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  pmos_prog.sym # of pins=8
** sym_path: /foss/designs/ttsky25a_minimosbius/xschem/pmos_prog.sym
** sch_path: /foss/designs/ttsky25a_minimosbius/xschem/pmos_prog.sch
.subckt pmos_prog VAPWR VDPWR Vs Vg Vd ctrl_source ctrl_width[1] ctrl_width[0] GND
*.ipin ctrl_width[1],ctrl_width[0]
*.iopin Vs
*.iopin Vg
*.iopin Vd
*.iopin VAPWR
*.iopin VDPWR
*.iopin GND
*.ipin ctrl_source
x1 GND VDPWR VAPWR ctrl_width[0] Vd_1x Vd tt_asw_3v3
x2 GND VDPWR VAPWR ctrl_width[1] Vd_2x Vd tt_asw_3v3
x3 GND VDPWR VAPWR ctrl_source Vs VAPWR tt_asw_3v3
XM1 Vd Vg Vs Vs sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=30 nf=6 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vd_1x Vg Vs Vs sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=30 nf=6 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vd_2x Vg Vs Vs sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=60 nf=12 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 Vs Vs Vs Vs sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 Vs Vs Vs Vs sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
