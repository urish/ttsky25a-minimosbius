magic
tech sky130A
magscale 1 2
timestamp 1757216467
<< dnwell >>
rect 8500 3200 10700 6700
rect 12200 3200 14400 6700
rect 38700 4500 42700 6750
rect 47100 4500 51100 6750
<< nwell >>
rect 8420 6494 10780 6780
rect 8420 3406 8706 6494
rect 10494 3406 10780 6494
rect 8420 3120 10780 3406
rect 12120 6494 14480 6780
rect 12120 3406 12406 6494
rect 14194 3406 14480 6494
rect 38620 6544 42780 6830
rect 38620 4706 38906 6544
rect 42494 4706 42780 6544
rect 38620 4420 42780 4706
rect 47020 6544 51180 6830
rect 47020 4706 47306 6544
rect 50894 4706 51180 6544
rect 47020 4420 51180 4706
rect 12120 3120 14480 3406
<< nsubdiff >>
rect 38657 6773 42743 6793
rect 8457 6723 10743 6743
rect 8457 6689 8537 6723
rect 10663 6689 10743 6723
rect 8457 6669 10743 6689
rect 8457 6663 8531 6669
rect 8457 3237 8477 6663
rect 8511 3237 8531 6663
rect 8457 3231 8531 3237
rect 10669 6663 10743 6669
rect 10669 3237 10689 6663
rect 10723 3237 10743 6663
rect 10669 3231 10743 3237
rect 8457 3211 10743 3231
rect 8457 3177 8537 3211
rect 10663 3177 10743 3211
rect 8457 3157 10743 3177
rect 12157 6723 14443 6743
rect 12157 6689 12237 6723
rect 14363 6689 14443 6723
rect 12157 6669 14443 6689
rect 12157 6663 12231 6669
rect 12157 3237 12177 6663
rect 12211 3237 12231 6663
rect 12157 3231 12231 3237
rect 14369 6663 14443 6669
rect 14369 3237 14389 6663
rect 14423 3237 14443 6663
rect 38657 6739 38737 6773
rect 42663 6739 42743 6773
rect 38657 6719 42743 6739
rect 38657 6713 38731 6719
rect 38657 4537 38677 6713
rect 38711 4537 38731 6713
rect 38657 4531 38731 4537
rect 42669 6713 42743 6719
rect 42669 4537 42689 6713
rect 42723 4537 42743 6713
rect 42669 4531 42743 4537
rect 38657 4511 42743 4531
rect 38657 4477 38737 4511
rect 42663 4477 42743 4511
rect 38657 4457 42743 4477
rect 47057 6773 51143 6793
rect 47057 6739 47137 6773
rect 51063 6739 51143 6773
rect 47057 6719 51143 6739
rect 47057 6713 47131 6719
rect 47057 4537 47077 6713
rect 47111 4537 47131 6713
rect 47057 4531 47131 4537
rect 51069 6713 51143 6719
rect 51069 4537 51089 6713
rect 51123 4537 51143 6713
rect 51069 4531 51143 4537
rect 47057 4511 51143 4531
rect 47057 4477 47137 4511
rect 51063 4477 51143 4511
rect 47057 4457 51143 4477
rect 14369 3231 14443 3237
rect 12157 3211 14443 3231
rect 12157 3177 12237 3211
rect 14363 3177 14443 3211
rect 12157 3157 14443 3177
<< nsubdiffcont >>
rect 8537 6689 10663 6723
rect 8477 3237 8511 6663
rect 10689 3237 10723 6663
rect 8537 3177 10663 3211
rect 12237 6689 14363 6723
rect 12177 3237 12211 6663
rect 14389 3237 14423 6663
rect 38737 6739 42663 6773
rect 38677 4537 38711 6713
rect 42689 4537 42723 6713
rect 38737 4477 42663 4511
rect 47137 6739 51063 6773
rect 47077 4537 47111 6713
rect 51089 4537 51123 6713
rect 47137 4477 51063 4511
rect 12237 3177 14363 3211
<< locali >>
rect 7900 7190 14900 7200
rect 7900 6710 8220 7190
rect 8900 6723 12010 7190
rect 12690 6723 14900 7190
rect 10663 6710 12010 6723
rect 7900 6689 8537 6710
rect 10663 6689 12237 6710
rect 14363 6689 14900 6723
rect 7900 6663 8511 6689
rect 7900 3237 8477 6663
rect 10689 6663 12211 6689
rect 8760 6260 10380 6460
rect 8760 6020 8960 6260
rect 10180 6040 10380 6260
rect 8760 5140 9100 6020
rect 10040 5160 10380 6040
rect 8760 4800 8960 5140
rect 10180 4800 10380 5160
rect 8760 3920 9100 4800
rect 10040 3920 10380 4800
rect 8760 3680 8960 3920
rect 10180 3680 10380 3920
rect 8760 3480 10380 3680
rect 7900 3211 8511 3237
rect 10723 3237 12177 6663
rect 14389 6663 14900 6689
rect 12460 6260 14080 6460
rect 12460 6020 12660 6260
rect 13880 6020 14080 6260
rect 12460 5140 12800 6020
rect 13740 5140 14080 6020
rect 12460 4800 12660 5140
rect 13880 4820 14080 5140
rect 12460 3920 12800 4800
rect 13740 3940 14080 4820
rect 12460 3680 12660 3920
rect 13880 3680 14080 3940
rect 12460 3480 14080 3680
rect 10689 3211 12211 3237
rect 14423 3237 14900 6663
rect 38290 6773 43100 7160
rect 38290 6739 38737 6773
rect 42663 6739 43100 6773
rect 38290 6713 38711 6739
rect 38290 5040 38677 6713
rect 42689 6713 43100 6739
rect 39030 6290 42320 6590
rect 39030 6100 39400 6290
rect 41950 6100 42320 6290
rect 39030 5120 39410 6100
rect 41930 5120 42320 6100
rect 38711 5040 38870 5050
rect 38290 4420 38630 5040
rect 38860 4511 38870 5040
rect 39030 4920 39400 5120
rect 41950 4920 42320 5120
rect 39030 4620 42320 4920
rect 42723 4537 43100 6713
rect 42689 4511 43100 4537
rect 42663 4477 43100 4511
rect 47077 6739 47137 6773
rect 51063 6739 51123 6773
rect 47077 6713 47111 6739
rect 51089 6713 51123 6739
rect 47430 6290 50720 6590
rect 47430 6100 47800 6290
rect 50350 6100 50720 6290
rect 47430 5120 47810 6100
rect 50330 5120 50720 6100
rect 47430 4920 47800 5120
rect 50350 4920 50720 5120
rect 47430 4620 50720 4920
rect 47077 4511 47111 4537
rect 51089 4511 51123 4537
rect 47077 4477 47137 4511
rect 51063 4477 51123 4511
rect 38860 4420 43100 4477
rect 38290 4100 43100 4420
rect 14389 3211 14900 3237
rect 7900 3177 8537 3211
rect 10663 3177 12237 3211
rect 14363 3177 14900 3211
rect 7900 2700 14900 3177
rect 38460 3470 46350 3670
rect 38460 3260 39000 3470
rect 45830 3260 46350 3470
rect 38460 2300 39070 3260
rect 45760 2300 46350 3260
rect 38460 2050 39000 2300
rect 38460 1090 39070 2050
rect 45830 2040 46350 2300
rect 38460 870 39000 1090
rect 45760 1080 46350 2040
rect 45840 870 46350 1080
rect 38460 670 46350 870
<< viali >>
rect 8220 6723 8900 7190
rect 12010 6723 12690 7190
rect 8220 6710 8537 6723
rect 8537 6710 8900 6723
rect 12010 6710 12237 6723
rect 12237 6710 12690 6723
rect 38630 4537 38677 5040
rect 38677 4537 38711 5040
rect 38711 4537 38860 5040
rect 38630 4511 38860 4537
rect 38630 4477 38737 4511
rect 38737 4477 38860 4511
rect 38630 4420 38860 4477
<< metal1 >>
rect 52930 9090 53290 9100
rect 52930 8490 53010 9090
rect 53280 8490 53290 9090
rect 52930 8480 53290 8490
rect 52930 7650 53230 8480
rect 8200 7190 8920 7200
rect 8200 6710 8220 7190
rect 8900 6710 8920 7190
rect 8200 6700 8920 6710
rect 11990 7190 12710 7200
rect 11990 6710 12010 7190
rect 12690 6710 12710 7190
rect 11990 6700 12710 6710
rect 13070 6200 13150 7580
rect 13390 6200 13470 7580
rect 52520 7400 53230 7650
rect 41180 7120 42520 7130
rect 41180 6840 41190 7120
rect 41560 6840 42210 7120
rect 42510 6840 42520 7120
rect 41180 6830 42520 6840
rect 39440 6410 45190 6420
rect 39440 6220 44800 6410
rect 8720 6120 10080 6200
rect 12780 6120 14100 6200
rect 8720 5040 8860 6120
rect 9880 6070 10040 6080
rect 9100 6060 9260 6070
rect 9100 5100 9110 6060
rect 9250 5100 9260 6060
rect 9100 5090 9260 5100
rect 9370 6060 9450 6070
rect 9370 5100 9380 6060
rect 9440 5100 9450 6060
rect 9370 5090 9450 5100
rect 9530 6060 9610 6070
rect 9530 5100 9540 6060
rect 9600 5100 9610 6060
rect 9530 5090 9610 5100
rect 9690 6060 9770 6070
rect 9690 5100 9700 6060
rect 9760 5100 9770 6060
rect 9880 5110 9890 6070
rect 10030 5110 10040 6070
rect 9880 5100 10040 5110
rect 12800 6060 12960 6070
rect 12800 5100 12810 6060
rect 12950 5100 12960 6060
rect 9690 5090 9770 5100
rect 12800 5090 12960 5100
rect 13070 6060 13150 6120
rect 13070 5100 13080 6060
rect 13140 5100 13150 6060
rect 13070 5090 13150 5100
rect 13230 6060 13310 6070
rect 13230 5100 13240 6060
rect 13300 5100 13310 6060
rect 13230 5090 13310 5100
rect 13390 6060 13470 6120
rect 13390 5100 13400 6060
rect 13460 5100 13470 6060
rect 13590 6060 13750 6070
rect 13590 6020 13600 6060
rect 13580 5140 13600 6020
rect 13390 5090 13470 5100
rect 13590 5100 13600 5140
rect 13740 5100 13750 6060
rect 13590 5090 13750 5100
rect 13960 5040 14100 6120
rect 39230 6100 39400 6190
rect 39460 6160 39510 6220
rect 39620 6160 39670 6220
rect 40090 6160 40140 6220
rect 40250 6160 40300 6220
rect 40720 6160 40770 6220
rect 40880 6160 40930 6220
rect 41350 6160 41400 6220
rect 41520 6160 41570 6220
rect 39230 6090 39420 6100
rect 39230 5130 39240 6090
rect 39410 5130 39420 6090
rect 39230 5120 39420 5130
rect 8720 4900 10080 5040
rect 12780 4900 14100 5040
rect 8720 4320 8860 4900
rect 8560 4310 8860 4320
rect 8560 4130 8570 4310
rect 8850 4130 8860 4310
rect 8560 4120 8860 4130
rect 8720 3820 8860 4120
rect 9100 4840 9260 4850
rect 9100 3880 9110 4840
rect 9250 3880 9260 4840
rect 9100 3870 9260 3880
rect 9370 4840 9450 4850
rect 9370 3880 9380 4840
rect 9440 3880 9450 4840
rect 9370 3870 9450 3880
rect 9530 4840 9610 4850
rect 9530 3880 9540 4840
rect 9600 3880 9610 4840
rect 9530 3870 9610 3880
rect 9690 4840 9770 4850
rect 9690 3880 9700 4840
rect 9760 3880 9770 4840
rect 9690 3870 9770 3880
rect 9880 4840 10040 4850
rect 9880 3880 9890 4840
rect 10030 3880 10040 4840
rect 9880 3870 10040 3880
rect 12800 4840 12960 4850
rect 12800 3880 12810 4840
rect 12950 3880 12960 4840
rect 12800 3870 12960 3880
rect 13070 4840 13150 4850
rect 13070 3880 13080 4840
rect 13140 3880 13150 4840
rect 13070 3870 13150 3880
rect 13230 4840 13310 4850
rect 13230 3880 13240 4840
rect 13300 3880 13310 4840
rect 13230 3870 13310 3880
rect 13390 4840 13470 4850
rect 13390 3880 13400 4840
rect 13460 3880 13470 4840
rect 13590 4840 13750 4850
rect 13590 4820 13600 4840
rect 13580 3940 13600 4820
rect 13390 3870 13470 3880
rect 13590 3880 13600 3940
rect 13740 3880 13750 4840
rect 13590 3870 13750 3880
rect 13960 4320 14100 4900
rect 38620 5040 38870 5060
rect 38620 4420 38630 5040
rect 38860 4420 38870 5040
rect 39230 5030 39400 5120
rect 39470 5050 39500 6160
rect 39540 6090 39600 6100
rect 39540 5120 39600 5130
rect 39630 5050 39660 6160
rect 39690 6090 39750 6100
rect 39690 5120 39750 5130
rect 39780 5050 39810 6160
rect 39850 6090 39910 6100
rect 39850 5120 39910 5130
rect 39940 5050 39970 6160
rect 40010 6090 40070 6100
rect 40010 5120 40070 5130
rect 40100 5050 40130 6160
rect 40170 6090 40230 6100
rect 40170 5120 40230 5130
rect 40260 5050 40290 6160
rect 40330 6090 40390 6100
rect 40330 5120 40390 5130
rect 40420 5050 40450 6160
rect 40480 6090 40540 6100
rect 40480 5120 40540 5130
rect 40580 5050 40610 6160
rect 40640 6090 40700 6100
rect 40640 5120 40700 5130
rect 40730 5050 40760 6160
rect 40800 6090 40860 6100
rect 40800 5120 40860 5130
rect 40890 5050 40920 6160
rect 40960 6090 41020 6100
rect 40960 5120 41020 5130
rect 41050 5050 41080 6160
rect 41120 6090 41180 6100
rect 41120 5120 41180 5130
rect 41210 5050 41240 6160
rect 41270 6090 41330 6100
rect 41270 5120 41330 5130
rect 41360 5050 41390 6160
rect 41430 6090 41490 6100
rect 41430 5120 41490 5130
rect 41530 5050 41560 6160
rect 41590 6090 41650 6100
rect 41590 5120 41650 5130
rect 41680 5050 41710 6160
rect 41750 6090 41810 6100
rect 41750 5120 41810 5130
rect 41850 5050 41880 6160
rect 41950 6100 42120 6190
rect 41930 6090 42120 6100
rect 41930 5130 41940 6090
rect 42110 5130 42120 6090
rect 44790 6030 44800 6220
rect 45180 6030 45190 6410
rect 47840 6410 51290 6420
rect 47840 6230 50730 6410
rect 51280 6230 51290 6410
rect 47840 6220 51290 6230
rect 44790 6020 45190 6030
rect 47560 6100 47800 6190
rect 47860 6160 47910 6220
rect 48020 6160 48070 6220
rect 48490 6160 48540 6220
rect 48650 6160 48700 6220
rect 49120 6160 49170 6220
rect 49280 6160 49330 6220
rect 49750 6160 49800 6220
rect 49920 6160 49970 6220
rect 47560 6090 47820 6100
rect 41930 5120 42120 5130
rect 39780 5000 39830 5050
rect 39930 5000 39980 5050
rect 40410 5000 40460 5050
rect 40570 5000 40620 5050
rect 41040 5000 41090 5050
rect 41200 5000 41250 5050
rect 41670 5000 41720 5050
rect 41840 5000 41890 5050
rect 41950 5030 42120 5120
rect 44190 5190 44590 5200
rect 44190 5000 44200 5190
rect 39440 4810 44200 5000
rect 44580 5000 44590 5190
rect 47560 5130 47640 6090
rect 47810 5130 47820 6090
rect 47560 5120 47820 5130
rect 44580 4810 45180 5000
rect 39440 4800 45180 4810
rect 38620 4400 38870 4420
rect 13960 4310 14260 4320
rect 13960 4130 13970 4310
rect 14250 4130 14260 4310
rect 47560 4290 47800 5120
rect 47870 5050 47900 6160
rect 47940 6090 48000 6100
rect 47940 5120 48000 5130
rect 48030 5050 48060 6160
rect 48090 6090 48150 6100
rect 48090 5120 48150 5130
rect 48180 5050 48210 6160
rect 48250 6090 48310 6100
rect 48250 5120 48310 5130
rect 48340 5050 48370 6160
rect 48410 6090 48470 6100
rect 48410 5120 48470 5130
rect 48500 5050 48530 6160
rect 48570 6090 48630 6100
rect 48570 5120 48630 5130
rect 48660 5050 48690 6160
rect 48730 6090 48790 6100
rect 48730 5120 48790 5130
rect 48820 5050 48850 6160
rect 48880 6090 48940 6100
rect 48880 5120 48940 5130
rect 48980 5050 49010 6160
rect 49040 6090 49100 6100
rect 49040 5120 49100 5130
rect 49130 5050 49160 6160
rect 49200 6090 49260 6100
rect 49200 5120 49260 5130
rect 49290 5050 49320 6160
rect 49360 6090 49420 6100
rect 49360 5120 49420 5130
rect 49450 5050 49480 6160
rect 49520 6090 49580 6100
rect 49520 5120 49580 5130
rect 49610 5050 49640 6160
rect 49670 6090 49730 6100
rect 49670 5120 49730 5130
rect 49760 5050 49790 6160
rect 49830 6090 49890 6100
rect 49830 5120 49890 5130
rect 49930 5050 49960 6160
rect 49990 6090 50050 6100
rect 49990 5120 50050 5130
rect 50080 5050 50110 6160
rect 50150 6090 50210 6100
rect 50150 5120 50210 5130
rect 50250 5050 50280 6160
rect 50350 6100 50520 6190
rect 50330 6090 50520 6100
rect 50330 5130 50340 6090
rect 50510 5800 50520 6090
rect 52520 5800 52920 7400
rect 50510 5400 52920 5800
rect 50510 5130 50520 5400
rect 50330 5120 50520 5130
rect 48180 5000 48230 5050
rect 48330 5000 48380 5050
rect 48810 5000 48860 5050
rect 48970 5000 49020 5050
rect 49440 5000 49490 5050
rect 49600 5000 49650 5050
rect 50070 5000 50120 5050
rect 50240 5000 50290 5050
rect 50350 5030 50520 5120
rect 52520 5330 52920 5400
rect 52520 5320 53300 5330
rect 47840 4990 51280 5000
rect 47840 4810 50720 4990
rect 51270 4810 51280 4990
rect 52520 4920 52530 5320
rect 53290 4920 53300 5320
rect 52520 4910 53300 4920
rect 47840 4800 51280 4810
rect 13960 4120 14260 4130
rect 47480 4280 47800 4290
rect 13960 3820 14100 4120
rect 47480 4100 47490 4280
rect 47790 4100 47800 4280
rect 47480 4090 47800 4100
rect 8720 3740 10080 3820
rect 12780 3740 14100 3820
rect 39080 3310 45720 3450
rect 38770 2700 39070 3270
rect 38770 2690 39090 2700
rect 38830 2310 39030 2690
rect 38770 2300 39090 2310
rect 38770 2040 39000 2300
rect 39150 2240 39230 3310
rect 39280 3250 39360 3260
rect 39280 2310 39290 3250
rect 39350 2310 39360 3250
rect 39280 2300 39360 2310
rect 39410 2240 39490 3310
rect 39540 2690 39600 2700
rect 39540 2300 39600 2310
rect 39660 2240 39740 3310
rect 39790 3250 39870 3260
rect 39790 2310 39800 3250
rect 39860 2310 39870 3250
rect 39790 2300 39870 2310
rect 39920 2240 40000 3310
rect 40060 2690 40120 2700
rect 40060 2300 40120 2310
rect 40180 2240 40260 3310
rect 40310 3240 40390 3260
rect 40310 2310 40320 3240
rect 40380 2310 40390 3240
rect 40310 2300 40390 2310
rect 40430 2240 40510 3310
rect 40580 2690 40640 2700
rect 40580 2300 40640 2310
rect 40700 2240 40780 3310
rect 40820 3250 40900 3260
rect 40820 2310 40830 3250
rect 40890 2310 40900 3250
rect 40820 2300 40900 2310
rect 40950 2240 41030 3310
rect 41090 2690 41150 2700
rect 41090 2300 41150 2310
rect 41210 2240 41290 3310
rect 41340 3250 41420 3260
rect 41340 2310 41350 3250
rect 41410 2310 41420 3250
rect 41340 2300 41420 2310
rect 41470 2240 41550 3310
rect 41610 2690 41670 2700
rect 41610 2300 41670 2310
rect 41730 2240 41810 3310
rect 41860 3250 41940 3260
rect 41860 2310 41870 3250
rect 41930 2310 41940 3250
rect 41860 2300 41940 2310
rect 41990 2240 42070 3310
rect 42120 2690 42180 2700
rect 42120 2300 42180 2310
rect 42250 2240 42330 3310
rect 42370 3250 42450 3260
rect 42370 2310 42380 3250
rect 42440 2310 42450 3250
rect 42370 2300 42450 2310
rect 42500 2240 42580 3310
rect 42640 2690 42700 2700
rect 42640 2300 42700 2310
rect 42760 2240 42840 3310
rect 42890 3250 42970 3260
rect 42890 2310 42900 3250
rect 42960 2310 42970 3250
rect 42890 2300 42970 2310
rect 43020 2240 43100 3310
rect 43160 2690 43220 2700
rect 43160 2300 43220 2310
rect 43280 2240 43360 3310
rect 43400 3250 43480 3260
rect 43400 2310 43410 3250
rect 43470 2310 43480 3250
rect 43400 2300 43480 2310
rect 43540 2240 43620 3310
rect 43670 2690 43730 2700
rect 43670 2300 43730 2310
rect 43790 2240 43870 3310
rect 43920 3250 44000 3260
rect 43920 2310 43930 3250
rect 43990 2310 44000 3250
rect 43920 2300 44000 2310
rect 44050 2240 44130 3310
rect 44190 2690 44250 2700
rect 44190 2300 44250 2310
rect 44310 2240 44390 3310
rect 44440 3250 44520 3260
rect 44440 2310 44450 3250
rect 44510 2310 44520 3250
rect 44440 2300 44520 2310
rect 44570 2240 44650 3310
rect 44700 2690 44760 2700
rect 44700 2300 44760 2310
rect 44820 2240 44900 3310
rect 44950 3250 45030 3260
rect 44950 2310 44960 3250
rect 45020 2310 45030 3250
rect 44950 2300 45030 2310
rect 45080 2240 45160 3310
rect 45220 2690 45280 2700
rect 45220 2300 45280 2310
rect 45340 2240 45420 3310
rect 45470 3250 45550 3260
rect 45470 2310 45480 3250
rect 45540 2310 45550 3250
rect 45470 2300 45550 2310
rect 45600 2240 45680 3310
rect 45750 2700 46040 3270
rect 45740 2690 46050 2700
rect 45800 2310 45990 2690
rect 45740 2300 45800 2310
rect 45830 2300 46050 2310
rect 39090 2230 45740 2240
rect 39090 2110 39100 2230
rect 39240 2110 39400 2230
rect 39750 2110 39910 2230
rect 40260 2110 40430 2230
rect 40780 2110 40940 2230
rect 41290 2110 41460 2230
rect 41810 2110 41980 2230
rect 42330 2110 42490 2230
rect 42840 2110 43010 2230
rect 43360 2110 43520 2230
rect 43870 2110 44040 2230
rect 44390 2110 44560 2230
rect 44910 2110 45070 2230
rect 45420 2110 45590 2230
rect 45730 2110 45740 2230
rect 39090 2100 45740 2110
rect 38770 1480 39080 2040
rect 38770 1470 39090 1480
rect 38830 1090 39030 1470
rect 38770 1080 39090 1090
rect 39150 1020 39230 2100
rect 39280 2030 39360 2040
rect 39280 1090 39290 2030
rect 39350 1090 39360 2030
rect 39280 1080 39360 1090
rect 39410 1020 39490 2100
rect 39540 1470 39600 1480
rect 39540 1080 39600 1090
rect 39660 1020 39740 2100
rect 39790 2030 39870 2040
rect 39790 1090 39800 2030
rect 39860 1090 39870 2030
rect 39790 1080 39870 1090
rect 39920 1020 40000 2100
rect 40060 1470 40120 1480
rect 40060 1080 40120 1090
rect 40180 1020 40260 2100
rect 40310 2030 40390 2040
rect 40310 1090 40320 2030
rect 40380 1090 40390 2030
rect 40310 1080 40390 1090
rect 40430 1020 40510 2100
rect 40580 1470 40640 1480
rect 40580 1080 40640 1090
rect 40700 1020 40780 2100
rect 40820 2030 40900 2040
rect 40820 1090 40830 2030
rect 40890 1090 40900 2030
rect 40820 1080 40900 1090
rect 40950 1020 41030 2100
rect 41090 1470 41150 1480
rect 41090 1080 41150 1090
rect 41210 1020 41550 2100
rect 41610 1470 41670 1480
rect 41610 1080 41670 1090
rect 41730 1020 41810 2100
rect 41860 2030 41940 2040
rect 41860 1090 41870 2030
rect 41930 1090 41940 2030
rect 41860 1080 41940 1090
rect 41990 1020 42070 2100
rect 42120 1470 42180 1480
rect 42120 1080 42180 1090
rect 42250 1020 42330 2100
rect 42370 2030 42450 2040
rect 42370 1090 42380 2030
rect 42440 1090 42450 2030
rect 42370 1080 42450 1090
rect 42500 1020 42580 2100
rect 42640 1470 42700 1480
rect 42640 1080 42700 1090
rect 42760 1020 42840 2100
rect 42890 2030 42970 2040
rect 42890 1090 42900 2030
rect 42960 1090 42970 2030
rect 42890 1080 42970 1090
rect 43020 1020 43100 2100
rect 43160 1470 43220 1480
rect 43160 1080 43220 1090
rect 43280 1020 43360 2100
rect 43400 2030 43480 2040
rect 43400 1090 43410 2030
rect 43470 1090 43480 2030
rect 43400 1080 43480 1090
rect 43540 1020 43620 2100
rect 43670 1470 43730 1480
rect 43670 1080 43730 1090
rect 43790 1020 43870 2100
rect 43920 2030 44000 2040
rect 43920 1090 43930 2030
rect 43990 1090 44000 2030
rect 43920 1080 44000 1090
rect 44050 1020 44130 2100
rect 44190 1470 44250 1480
rect 44190 1080 44250 1090
rect 44310 1020 44390 2100
rect 44440 2030 44520 2040
rect 44440 1090 44450 2030
rect 44510 1090 44520 2030
rect 44440 1080 44520 1090
rect 44570 1020 44650 2100
rect 44700 1470 44760 1480
rect 44700 1080 44760 1090
rect 44820 1020 44900 2100
rect 44950 2030 45030 2040
rect 44950 1090 44960 2030
rect 45020 1090 45030 2030
rect 44950 1080 45030 1090
rect 45080 1020 45160 2100
rect 45220 1470 45280 1480
rect 45220 1080 45280 1090
rect 45340 1020 45420 2100
rect 45470 2030 45550 2040
rect 45470 1090 45480 2030
rect 45540 1090 45550 2030
rect 45470 1080 45550 1090
rect 45600 1020 45680 2100
rect 45830 2040 46040 2300
rect 45750 1480 46040 2040
rect 45740 1470 46050 1480
rect 45800 1090 45990 1470
rect 45740 1080 46050 1090
rect 39090 880 45730 1020
<< via1 >>
rect 53010 8490 53280 9090
rect 8220 6710 8900 7190
rect 12010 6710 12690 7190
rect 41190 6840 41560 7120
rect 42210 6840 42510 7120
rect 9110 5100 9250 6060
rect 9380 5100 9440 6060
rect 9540 5100 9600 6060
rect 9700 5100 9760 6060
rect 9890 5110 10030 6070
rect 12810 5100 12950 6060
rect 13080 5100 13140 6060
rect 13240 5100 13300 6060
rect 13400 5100 13460 6060
rect 13600 5100 13740 6060
rect 39240 5130 39410 6090
rect 8570 4130 8850 4310
rect 9110 3880 9250 4840
rect 9380 3880 9440 4840
rect 9540 3880 9600 4840
rect 9700 3880 9760 4840
rect 9890 3880 10030 4840
rect 12810 3880 12950 4840
rect 13080 3880 13140 4840
rect 13240 3880 13300 4840
rect 13400 3880 13460 4840
rect 13600 3880 13740 4840
rect 38630 4420 38860 5040
rect 39540 5130 39600 6090
rect 39690 5130 39750 6090
rect 39850 5130 39910 6090
rect 40010 5130 40070 6090
rect 40170 5130 40230 6090
rect 40330 5130 40390 6090
rect 40480 5130 40540 6090
rect 40640 5130 40700 6090
rect 40800 5130 40860 6090
rect 40960 5130 41020 6090
rect 41120 5130 41180 6090
rect 41270 5130 41330 6090
rect 41430 5130 41490 6090
rect 41590 5130 41650 6090
rect 41750 5130 41810 6090
rect 41940 5130 42110 6090
rect 44800 6030 45180 6410
rect 50730 6230 51280 6410
rect 44200 4810 44580 5190
rect 47640 5130 47810 6090
rect 13970 4130 14250 4310
rect 47940 5130 48000 6090
rect 48090 5130 48150 6090
rect 48250 5130 48310 6090
rect 48410 5130 48470 6090
rect 48570 5130 48630 6090
rect 48730 5130 48790 6090
rect 48880 5130 48940 6090
rect 49040 5130 49100 6090
rect 49200 5130 49260 6090
rect 49360 5130 49420 6090
rect 49520 5130 49580 6090
rect 49670 5130 49730 6090
rect 49830 5130 49890 6090
rect 49990 5130 50050 6090
rect 50150 5130 50210 6090
rect 50340 5130 50510 6090
rect 50720 4810 51270 4990
rect 52530 4920 53290 5320
rect 47490 4100 47790 4280
rect 38770 2310 38830 2690
rect 39030 2310 39090 2690
rect 39290 2310 39350 3250
rect 39540 2310 39600 2690
rect 39800 2310 39860 3250
rect 40060 2310 40120 2690
rect 40320 2310 40380 3240
rect 40580 2310 40640 2690
rect 40830 2310 40890 3250
rect 41090 2310 41150 2690
rect 41350 2310 41410 3250
rect 41610 2310 41670 2690
rect 41870 2310 41930 3250
rect 42120 2310 42180 2690
rect 42380 2310 42440 3250
rect 42640 2310 42700 2690
rect 42900 2310 42960 3250
rect 43160 2310 43220 2690
rect 43410 2310 43470 3250
rect 43670 2310 43730 2690
rect 43930 2310 43990 3250
rect 44190 2310 44250 2690
rect 44450 2310 44510 3250
rect 44700 2310 44760 2690
rect 44960 2310 45020 3250
rect 45220 2310 45280 2690
rect 45480 2310 45540 3250
rect 45740 2310 45800 2690
rect 45990 2310 46050 2690
rect 39100 2110 39240 2230
rect 39400 2110 39750 2230
rect 39910 2110 40260 2230
rect 40430 2110 40780 2230
rect 40940 2110 41290 2230
rect 41460 2110 41810 2230
rect 41980 2110 42330 2230
rect 42490 2110 42840 2230
rect 43010 2110 43360 2230
rect 43520 2110 43870 2230
rect 44040 2110 44390 2230
rect 44560 2110 44910 2230
rect 45070 2110 45420 2230
rect 45590 2110 45730 2230
rect 38770 1090 38830 1470
rect 39030 1090 39090 1470
rect 39290 1090 39350 2030
rect 39540 1090 39600 1470
rect 39800 1090 39860 2030
rect 40060 1090 40120 1470
rect 40320 1090 40380 2030
rect 40580 1090 40640 1470
rect 40830 1090 40890 2030
rect 41090 1090 41150 1470
rect 41610 1090 41670 1470
rect 41870 1090 41930 2030
rect 42120 1090 42180 1470
rect 42380 1090 42440 2030
rect 42640 1090 42700 1470
rect 42900 1090 42960 2030
rect 43160 1090 43220 1470
rect 43410 1090 43470 2030
rect 43670 1090 43730 1470
rect 43930 1090 43990 2030
rect 44190 1090 44250 1470
rect 44450 1090 44510 2030
rect 44700 1090 44760 1470
rect 44960 1090 45020 2030
rect 45220 1090 45280 1470
rect 45480 1090 45540 2030
rect 45740 1090 45800 1470
rect 45990 1090 46050 1470
<< metal2 >>
rect 53000 9090 53290 9100
rect 15740 8330 16400 8340
rect 3380 8250 3860 8260
rect 3380 7710 3390 8250
rect 3850 7710 3860 8250
rect 15740 7970 15750 8330
rect 16390 7970 16400 8330
rect 15740 7960 16400 7970
rect 19510 8320 19990 8330
rect 12950 7900 13220 7910
rect 3380 7700 3860 7710
rect 9250 7890 9520 7900
rect 9250 7580 9260 7890
rect 9510 7580 9520 7890
rect 9250 7570 9520 7580
rect 9620 7890 9890 7900
rect 9620 7580 9630 7890
rect 9880 7580 9890 7890
rect 12950 7590 12960 7900
rect 13210 7590 13220 7900
rect 12950 7580 13220 7590
rect 13320 7900 13590 7910
rect 13320 7590 13330 7900
rect 13580 7590 13590 7900
rect 19510 7780 19520 8320
rect 19980 7780 19990 8320
rect 19510 7770 19990 7780
rect 13320 7580 13590 7590
rect 9620 7570 9890 7580
rect 8200 7190 8920 7200
rect 8200 6710 8220 7190
rect 8900 6710 8920 7190
rect 8200 6700 8920 6710
rect 9100 6060 9260 6070
rect 9100 5100 9110 6060
rect 9250 5100 9260 6060
rect 9100 5090 9260 5100
rect 9370 6060 9450 7570
rect 9370 5100 9380 6060
rect 9440 5100 9450 6060
rect 9370 5090 9450 5100
rect 9530 6060 9610 6070
rect 9530 5100 9540 6060
rect 9600 5100 9610 6060
rect 9530 5090 9610 5100
rect 9690 6060 9770 7570
rect 12000 7190 12700 7200
rect 12000 6710 12010 7190
rect 12690 6710 12700 7190
rect 12000 6700 12700 6710
rect 9690 5100 9700 6060
rect 9760 5100 9770 6060
rect 9880 6070 10040 6080
rect 9880 5110 9890 6070
rect 10030 5110 10040 6070
rect 9880 5100 10040 5110
rect 12800 6060 12960 6070
rect 12800 5100 12810 6060
rect 12950 5100 12960 6060
rect 9100 4840 9260 4850
rect 8560 4310 8860 4320
rect 8560 4130 8570 4310
rect 8850 4130 8860 4310
rect 8560 4120 8860 4130
rect 9100 3880 9110 4840
rect 9250 3880 9260 4840
rect 9100 3870 9260 3880
rect 9370 4840 9450 4850
rect 9370 3880 9380 4840
rect 9440 3880 9450 4840
rect 9370 3870 9450 3880
rect 9530 4840 9610 4850
rect 9530 3880 9540 4840
rect 9600 3880 9610 4840
rect 9530 3870 9610 3880
rect 9690 4840 9770 5100
rect 12800 5090 12960 5100
rect 13070 6060 13150 7580
rect 13070 5100 13080 6060
rect 13140 5100 13150 6060
rect 9690 3880 9700 4840
rect 9760 3880 9770 4840
rect 9690 3870 9770 3880
rect 9880 4840 10040 4850
rect 9880 3880 9890 4840
rect 10030 3880 10040 4840
rect 9880 3870 10040 3880
rect 12800 4840 12960 4850
rect 12800 3880 12810 4840
rect 12950 3880 12960 4840
rect 12800 3870 12960 3880
rect 13070 4840 13150 5100
rect 13230 6060 13310 6070
rect 13230 5100 13240 6060
rect 13300 5100 13310 6060
rect 13230 5090 13310 5100
rect 13390 6060 13470 7580
rect 13390 5100 13400 6060
rect 13460 5100 13470 6060
rect 13390 5090 13470 5100
rect 13590 6060 13750 6070
rect 13590 5100 13600 6060
rect 13740 5100 13750 6060
rect 37970 5800 38250 8620
rect 41180 7120 41570 8560
rect 41180 6840 41190 7120
rect 41560 6840 41570 7120
rect 41180 6830 41570 6840
rect 41740 6700 42030 8880
rect 53000 8490 53010 9090
rect 53280 8490 53290 9090
rect 53000 8480 53290 8490
rect 42200 7120 42520 7130
rect 42200 6840 42210 7120
rect 42510 6840 42520 7120
rect 42200 6830 42520 6840
rect 41740 6520 42130 6700
rect 39440 6450 41660 6460
rect 39440 6270 39450 6450
rect 41650 6270 41660 6450
rect 39440 6260 41660 6270
rect 39230 6090 39420 6100
rect 37950 5790 38280 5800
rect 37950 5410 37960 5790
rect 38270 5410 38280 5790
rect 37950 5400 38280 5410
rect 39230 5130 39240 6090
rect 39410 5130 39420 6090
rect 39230 5120 39420 5130
rect 39530 6090 39610 6260
rect 39530 5130 39540 6090
rect 39600 5130 39610 6090
rect 39530 5120 39610 5130
rect 39680 6090 39760 6100
rect 39680 5130 39690 6090
rect 39750 5130 39760 6090
rect 39680 5120 39760 5130
rect 39840 6090 39920 6100
rect 39840 5130 39850 6090
rect 39910 5130 39920 6090
rect 13590 5090 13750 5100
rect 38620 5040 38870 5050
rect 13070 3880 13080 4840
rect 13140 3880 13150 4840
rect 13070 3870 13150 3880
rect 13230 4840 13310 4850
rect 13230 3880 13240 4840
rect 13300 3880 13310 4840
rect 13230 3870 13310 3880
rect 13390 4840 13470 4850
rect 13390 3810 13400 4840
rect 13460 3810 13470 4840
rect 13590 4840 13750 4850
rect 13590 3880 13600 4840
rect 13740 3880 13750 4840
rect 38620 4420 38630 5040
rect 38860 4420 38870 5040
rect 39840 4950 39920 5130
rect 40000 6090 40080 6100
rect 40000 5130 40010 6090
rect 40070 5130 40080 6090
rect 40000 5120 40080 5130
rect 40160 6090 40240 6260
rect 40160 5130 40170 6090
rect 40230 5130 40240 6090
rect 40160 5120 40240 5130
rect 40320 6090 40400 6100
rect 40320 5130 40330 6090
rect 40390 5130 40400 6090
rect 40320 5120 40400 5130
rect 40470 6090 40550 6100
rect 40470 5130 40480 6090
rect 40540 5130 40550 6090
rect 40470 4950 40550 5130
rect 40630 6090 40710 6100
rect 40630 5130 40640 6090
rect 40700 5130 40710 6090
rect 40630 5120 40710 5130
rect 40790 6090 40870 6260
rect 40790 5130 40800 6090
rect 40860 5130 40870 6090
rect 40790 5120 40870 5130
rect 40950 6090 41030 6100
rect 40950 5130 40960 6090
rect 41020 5130 41030 6090
rect 40950 5120 41030 5130
rect 41110 6090 41190 6100
rect 41110 5130 41120 6090
rect 41180 5130 41190 6090
rect 41110 4950 41190 5130
rect 41260 6090 41340 6100
rect 41260 5130 41270 6090
rect 41330 5130 41340 6090
rect 41260 5120 41340 5130
rect 41420 6090 41500 6260
rect 41420 5130 41430 6090
rect 41490 5130 41500 6090
rect 41420 5120 41500 5130
rect 41580 6090 41660 6100
rect 41580 5130 41590 6090
rect 41650 5130 41660 6090
rect 41580 5120 41660 5130
rect 41740 6090 41820 6100
rect 41740 5130 41750 6090
rect 41810 5130 41820 6090
rect 41740 4950 41820 5130
rect 39440 4940 41820 4950
rect 39440 4760 39450 4940
rect 41810 4760 41820 4940
rect 39440 4750 41820 4760
rect 41930 6090 42130 6520
rect 41930 5130 41940 6090
rect 42110 5130 42130 6090
rect 38620 4410 38870 4420
rect 13960 4310 14260 4320
rect 13960 4130 13970 4310
rect 14250 4130 14260 4310
rect 40760 4250 40960 4260
rect 13960 4120 14260 4130
rect 13590 3870 13750 3880
rect 13390 3800 13470 3810
rect 33640 960 34020 4200
rect 40760 3870 40770 4250
rect 40950 3870 40960 4250
rect 41930 3900 42130 5130
rect 40760 3860 40960 3870
rect 37410 3260 37800 3840
rect 39730 3720 39930 3730
rect 39730 3340 39740 3720
rect 39920 3340 39930 3720
rect 39730 3330 39930 3340
rect 37410 3250 39360 3260
rect 37410 2840 39290 3250
rect 38770 2690 38830 2700
rect 38770 2300 38830 2310
rect 39030 2690 39090 2700
rect 39030 2300 39090 2310
rect 39280 2310 39290 2840
rect 39350 2310 39360 3250
rect 39790 3250 39870 3330
rect 39280 2300 39360 2310
rect 39540 2690 39600 2700
rect 39540 2300 39600 2310
rect 39790 2310 39800 3250
rect 39860 2310 39870 3250
rect 40820 3250 40900 3860
rect 40250 3230 40320 3240
rect 40380 3230 40450 3240
rect 40250 2850 40260 3230
rect 40440 2850 40450 3230
rect 40250 2840 40320 2850
rect 39790 2300 39870 2310
rect 40060 2690 40120 2700
rect 40060 2300 40120 2310
rect 40310 2310 40320 2840
rect 40380 2840 40450 2850
rect 40380 2310 40390 2840
rect 39090 2230 39250 2240
rect 39090 2110 39100 2230
rect 39240 2110 39250 2230
rect 39090 2100 39250 2110
rect 39390 2230 39760 2240
rect 39390 2110 39400 2230
rect 39750 2110 39760 2230
rect 39390 2100 39760 2110
rect 39900 2230 40270 2240
rect 39900 2110 39910 2230
rect 40260 2110 40270 2230
rect 39900 2100 40270 2110
rect 39280 2030 39360 2040
rect 39280 2000 39290 2030
rect 39220 1990 39290 2000
rect 39350 2000 39360 2030
rect 39790 2030 39870 2040
rect 39350 1990 39420 2000
rect 39220 1610 39230 1990
rect 39410 1610 39420 1990
rect 39220 1600 39290 1610
rect 38770 1470 38830 1480
rect 38770 1080 38830 1090
rect 39030 1470 39090 1480
rect 39030 1080 39090 1090
rect 39280 1090 39290 1600
rect 39350 1600 39420 1610
rect 39350 1090 39360 1600
rect 39280 1080 39360 1090
rect 39540 1470 39600 1480
rect 39540 1080 39600 1090
rect 39790 1090 39800 2030
rect 39860 1090 39870 2030
rect 40310 2030 40390 2310
rect 40580 2690 40640 2700
rect 40580 2300 40640 2310
rect 40820 2310 40830 3250
rect 40890 2310 40900 3250
rect 41340 3690 42130 3900
rect 41340 3250 41420 3690
rect 40420 2230 40790 2240
rect 40420 2110 40430 2230
rect 40780 2110 40790 2230
rect 40420 2100 40790 2110
rect 39790 970 39870 1090
rect 40060 1470 40120 1480
rect 40060 1080 40120 1090
rect 40310 1090 40320 2030
rect 40380 1090 40390 2030
rect 40820 2030 40900 2310
rect 41090 2690 41150 2700
rect 41090 2300 41150 2310
rect 41340 2310 41350 3250
rect 41410 2310 41420 3250
rect 41860 3250 41940 3690
rect 42320 3260 42520 6830
rect 42830 3740 43030 8030
rect 44790 6410 45190 6420
rect 44790 6030 44800 6410
rect 45180 6030 45190 6410
rect 44790 6020 45190 6030
rect 45530 5790 45930 8350
rect 53450 7760 53840 8340
rect 51920 7470 53840 7760
rect 47840 6450 50060 6460
rect 47840 6270 47850 6450
rect 50050 6270 50060 6450
rect 47840 6260 50060 6270
rect 50720 6410 51290 6420
rect 45530 5410 45540 5790
rect 45920 5410 45930 5790
rect 45530 5400 45930 5410
rect 47630 6090 47820 6100
rect 44190 5190 44590 5200
rect 44190 4810 44200 5190
rect 44580 4810 44590 5190
rect 47630 5130 47640 6090
rect 47810 5130 47820 6090
rect 47630 5120 47820 5130
rect 47930 6090 48010 6260
rect 47930 5130 47940 6090
rect 48000 5130 48010 6090
rect 47930 5120 48010 5130
rect 48080 6090 48160 6100
rect 48080 5130 48090 6090
rect 48150 5130 48160 6090
rect 48080 5120 48160 5130
rect 48240 6090 48320 6100
rect 48240 5130 48250 6090
rect 48310 5130 48320 6090
rect 48240 4950 48320 5130
rect 48400 6090 48480 6100
rect 48400 5130 48410 6090
rect 48470 5130 48480 6090
rect 48400 5120 48480 5130
rect 48560 6090 48640 6260
rect 48560 5130 48570 6090
rect 48630 5130 48640 6090
rect 48560 5120 48640 5130
rect 48720 6090 48800 6100
rect 48720 5130 48730 6090
rect 48790 5130 48800 6090
rect 48720 5120 48800 5130
rect 48870 6090 48950 6100
rect 48870 5130 48880 6090
rect 48940 5130 48950 6090
rect 48870 4950 48950 5130
rect 49030 6090 49110 6100
rect 49030 5130 49040 6090
rect 49100 5130 49110 6090
rect 49030 5120 49110 5130
rect 49190 6090 49270 6260
rect 49190 5130 49200 6090
rect 49260 5130 49270 6090
rect 49190 5120 49270 5130
rect 49350 6090 49430 6100
rect 49350 5130 49360 6090
rect 49420 5130 49430 6090
rect 49350 5120 49430 5130
rect 49510 6090 49590 6100
rect 49510 5130 49520 6090
rect 49580 5130 49590 6090
rect 49510 4950 49590 5130
rect 49660 6090 49740 6100
rect 49660 5130 49670 6090
rect 49730 5130 49740 6090
rect 49660 5120 49740 5130
rect 49820 6090 49900 6260
rect 50720 6230 50730 6410
rect 51280 6230 51290 6410
rect 50720 6220 51290 6230
rect 49820 5130 49830 6090
rect 49890 5130 49900 6090
rect 49820 5120 49900 5130
rect 49980 6090 50060 6100
rect 49980 5130 49990 6090
rect 50050 5130 50060 6090
rect 49980 5120 50060 5130
rect 50140 6090 50220 6100
rect 50140 5130 50150 6090
rect 50210 5130 50220 6090
rect 50140 4950 50220 5130
rect 50330 6090 50530 6100
rect 50330 5130 50340 6090
rect 50510 5130 50530 6090
rect 50330 5120 50530 5130
rect 44190 4800 44590 4810
rect 47840 4940 50220 4950
rect 47840 4760 47850 4940
rect 50210 4760 50220 4940
rect 50710 4990 51280 5000
rect 50710 4810 50720 4990
rect 51270 4810 51280 4990
rect 50710 4800 51280 4810
rect 47840 4750 50220 4760
rect 43860 4280 44590 4290
rect 43860 4100 43870 4280
rect 44580 4100 44590 4280
rect 43860 4090 44590 4100
rect 47480 4280 47800 4290
rect 47480 4100 47490 4280
rect 47790 4100 47800 4280
rect 47480 4090 47800 4100
rect 51920 4230 52310 7470
rect 52520 5320 53300 5330
rect 52520 4920 52530 5320
rect 53290 4920 53300 5320
rect 52520 4910 53300 4920
rect 42830 3540 43550 3740
rect 42830 3260 43030 3540
rect 41340 2300 41420 2310
rect 41610 2690 41670 2700
rect 41610 2300 41670 2310
rect 41860 2310 41870 3250
rect 41930 2310 41940 3250
rect 42370 3250 42450 3260
rect 41860 2300 41940 2310
rect 42120 2690 42180 2700
rect 42120 2300 42180 2310
rect 42370 2310 42380 3250
rect 42440 2310 42450 3250
rect 42890 3250 42970 3260
rect 43350 3250 43550 3540
rect 43860 3260 44060 4090
rect 44380 4010 45110 4020
rect 44380 3830 44390 4010
rect 45100 3830 45110 4010
rect 44380 3820 45110 3830
rect 51920 3830 51930 4230
rect 52300 3830 52310 4230
rect 51920 3820 52310 3830
rect 44380 3260 44580 3820
rect 44890 3740 45620 3750
rect 44890 3560 44900 3740
rect 45610 3560 45620 3740
rect 44890 3550 45620 3560
rect 44890 3260 45090 3550
rect 45410 3260 45610 3550
rect 43920 3250 44000 3260
rect 40930 2230 41300 2240
rect 40930 2110 40940 2230
rect 41290 2110 41300 2230
rect 40930 2100 41300 2110
rect 41450 2230 41820 2240
rect 41450 2110 41460 2230
rect 41810 2110 41820 2230
rect 41450 2100 41820 2110
rect 41970 2230 42340 2240
rect 41970 2110 41980 2230
rect 42330 2110 42340 2230
rect 41970 2100 42340 2110
rect 40310 1080 40390 1090
rect 40580 1470 40640 1480
rect 40580 1080 40640 1090
rect 40820 1090 40830 2030
rect 40890 1090 40900 2030
rect 41860 2030 41940 2040
rect 40820 1080 40900 1090
rect 41090 1470 41150 1480
rect 41090 1080 41150 1090
rect 41610 1470 41670 1480
rect 41610 1080 41670 1090
rect 41860 1090 41870 2030
rect 41930 1090 41940 2030
rect 42370 2030 42450 2310
rect 42640 2690 42700 2700
rect 42640 2300 42700 2310
rect 42890 2310 42900 3250
rect 42960 2310 42970 3250
rect 42480 2230 42850 2240
rect 42480 2110 42490 2230
rect 42840 2110 42850 2230
rect 42480 2100 42850 2110
rect 33640 580 33650 960
rect 34010 580 34020 960
rect 33640 570 34020 580
rect 39730 960 39930 970
rect 39730 580 39740 960
rect 39920 580 39930 960
rect 41860 740 41940 1090
rect 42120 1470 42180 1480
rect 42120 1080 42180 1090
rect 42370 1090 42380 2030
rect 42440 1090 42450 2030
rect 42890 2030 42970 2310
rect 43160 2690 43220 2700
rect 43160 2300 43220 2310
rect 43400 2310 43410 3250
rect 43470 2310 43480 3250
rect 43000 2230 43370 2240
rect 43000 2110 43010 2230
rect 43360 2110 43370 2230
rect 43000 2100 43370 2110
rect 42370 1080 42450 1090
rect 42640 1470 42700 1480
rect 42640 1080 42700 1090
rect 42890 1090 42900 2030
rect 42960 1090 42970 2030
rect 43400 2030 43480 2310
rect 43670 2690 43730 2700
rect 43670 2300 43730 2310
rect 43920 2310 43930 3250
rect 43990 2310 44000 3250
rect 44440 3250 44520 3260
rect 43510 2230 43880 2240
rect 43510 2110 43520 2230
rect 43870 2110 43880 2230
rect 43510 2100 43880 2110
rect 42890 1080 42970 1090
rect 43160 1470 43220 1480
rect 43160 1080 43220 1090
rect 43400 1090 43410 2030
rect 43470 1090 43480 2030
rect 43920 2030 44000 2310
rect 44190 2690 44250 2700
rect 44190 2300 44250 2310
rect 44440 2310 44450 3250
rect 44510 2310 44520 3250
rect 44950 3250 45030 3260
rect 44030 2230 44400 2240
rect 44030 2110 44040 2230
rect 44390 2110 44400 2230
rect 44030 2100 44400 2110
rect 43400 1080 43480 1090
rect 43670 1470 43730 1480
rect 43670 1080 43730 1090
rect 43920 1090 43930 2030
rect 43990 1090 44000 2030
rect 44440 2030 44520 2310
rect 44700 2690 44760 2700
rect 44700 2300 44760 2310
rect 44950 2310 44960 3250
rect 45020 2310 45030 3250
rect 45470 3250 45550 3260
rect 44550 2230 44920 2240
rect 44550 2110 44560 2230
rect 44910 2110 44920 2230
rect 44550 2100 44920 2110
rect 43920 1080 44000 1090
rect 44190 1470 44250 1480
rect 44190 1080 44250 1090
rect 44440 1090 44450 2030
rect 44510 1090 44520 2030
rect 44950 2030 45030 2310
rect 45220 2690 45280 2700
rect 45220 2300 45280 2310
rect 45470 2310 45480 3250
rect 45540 2310 45550 3250
rect 45060 2230 45430 2240
rect 45060 2110 45070 2230
rect 45420 2110 45430 2230
rect 45060 2100 45430 2110
rect 44440 1080 44520 1090
rect 44700 1470 44760 1480
rect 44700 1080 44760 1090
rect 44950 1090 44960 2030
rect 45020 1090 45030 2030
rect 45470 2030 45550 2310
rect 45740 2690 45800 2700
rect 45740 2300 45800 2310
rect 45990 2690 46050 2700
rect 45990 2300 46050 2310
rect 45580 2230 45740 2240
rect 45580 2110 45590 2230
rect 45730 2110 45740 2230
rect 45580 2100 45740 2110
rect 44950 1080 45030 1090
rect 45220 1470 45280 1480
rect 45220 1080 45280 1090
rect 45470 1090 45480 2030
rect 45540 1090 45550 2030
rect 45470 1080 45550 1090
rect 45740 1470 45800 1480
rect 45740 1080 45800 1090
rect 45990 1470 46050 1480
rect 45990 1080 46050 1090
rect 39730 570 39930 580
<< via2 >>
rect 3390 7710 3850 8250
rect 6970 7970 7610 8330
rect 15750 7970 16390 8330
rect 9260 7580 9510 7890
rect 9630 7580 9880 7890
rect 12960 7590 13210 7900
rect 13330 7590 13580 7900
rect 19520 7780 19980 8320
rect 8220 6710 8900 7190
rect 9110 5140 9250 5440
rect 9540 5140 9600 5440
rect 12010 6710 12690 7190
rect 9890 5140 10030 5440
rect 12810 5140 12950 5440
rect 8570 4130 8850 4310
rect 9110 4500 9250 4800
rect 9380 3880 9440 4480
rect 9540 4500 9600 4800
rect 9890 4500 10030 4800
rect 12810 4500 12950 4800
rect 13240 5140 13300 5440
rect 13600 5140 13740 5440
rect 39450 6270 41650 6450
rect 37960 5410 38270 5790
rect 39240 5410 39410 5790
rect 39690 5410 39750 5790
rect 13240 4500 13300 4800
rect 13400 3880 13460 4480
rect 13400 3810 13460 3880
rect 13600 4500 13740 4800
rect 38630 4420 38860 5040
rect 40010 5410 40070 5790
rect 40330 5410 40390 5790
rect 40640 5410 40700 5790
rect 40960 5410 41020 5790
rect 41270 5410 41330 5790
rect 41590 5410 41650 5790
rect 39450 4760 41810 4940
rect 41940 5410 42110 5790
rect 13970 4130 14250 4310
rect 40770 3870 40950 4250
rect 39740 3340 39920 3720
rect 38770 2310 38830 2690
rect 39030 2310 39090 2690
rect 39540 2310 39600 2690
rect 40260 2850 40320 3230
rect 40320 2850 40380 3230
rect 40380 2850 40440 3230
rect 40060 2310 40120 2690
rect 39100 2110 39240 2230
rect 39400 2110 39750 2230
rect 39910 2110 40260 2230
rect 39230 1610 39290 1990
rect 39290 1610 39350 1990
rect 39350 1610 39410 1990
rect 38770 1090 38830 1470
rect 39030 1090 39090 1470
rect 39540 1090 39600 1470
rect 40580 2310 40640 2690
rect 40430 2110 40780 2230
rect 40060 1090 40120 1470
rect 41090 2310 41150 2690
rect 44800 6030 45180 6410
rect 47850 6270 50050 6450
rect 45540 5410 45920 5790
rect 44200 4810 44580 5190
rect 47640 5410 47810 5790
rect 48090 5410 48150 5790
rect 48410 5410 48470 5790
rect 48730 5410 48790 5790
rect 49040 5410 49100 5790
rect 49360 5410 49420 5790
rect 49670 5410 49730 5790
rect 50730 6230 51280 6410
rect 49990 5410 50050 5790
rect 50340 5410 50510 5790
rect 47850 4760 50210 4940
rect 50720 4810 51270 4990
rect 43870 4100 44580 4280
rect 47490 4100 47790 4280
rect 41610 2310 41670 2690
rect 42120 2310 42180 2690
rect 44390 3830 45100 4010
rect 51930 3830 52300 4230
rect 44900 3560 45610 3740
rect 56280 3340 56650 3740
rect 40940 2110 41290 2230
rect 41460 2110 41810 2230
rect 41980 2110 42330 2230
rect 40580 1090 40640 1470
rect 41090 1090 41150 1470
rect 41610 1090 41670 1470
rect 42640 2310 42700 2690
rect 42490 2110 42840 2230
rect 33650 580 34010 960
rect 39740 580 39920 960
rect 42120 1090 42180 1470
rect 43160 2310 43220 2690
rect 43010 2110 43360 2230
rect 42640 1090 42700 1470
rect 43670 2310 43730 2690
rect 43520 2110 43870 2230
rect 43160 1090 43220 1470
rect 44190 2310 44250 2690
rect 44040 2110 44390 2230
rect 43670 1090 43730 1470
rect 44700 2310 44760 2690
rect 44560 2110 44910 2230
rect 44190 1090 44250 1470
rect 45220 2310 45280 2690
rect 45070 2110 45420 2230
rect 44700 1090 44760 1470
rect 45740 2310 45800 2690
rect 45990 2310 46050 2690
rect 45590 2110 45730 2230
rect 45220 1090 45280 1470
rect 45740 1090 45800 1470
rect 45990 1090 46050 1470
<< metal3 >>
rect 27310 39380 27550 39390
rect 23220 39370 24260 39380
rect 23450 39190 24260 39370
rect 23220 38990 24260 39190
rect 27310 38760 27320 39380
rect 27540 38990 28140 39380
rect 27540 38760 27550 38990
rect 27310 38560 27550 38760
rect 1880 36800 2280 37660
rect 5652 36800 6052 37300
rect 9424 36800 9824 37300
rect 24512 36800 24912 37300
rect 28284 36800 28684 37300
rect 32056 36800 32456 37300
rect 39600 36800 40000 37300
rect 43372 36800 43772 37300
rect 50916 36800 51316 37300
rect 54688 36800 55088 37300
rect 58460 36800 58860 37300
rect 69776 36800 70176 37300
rect 73548 36800 73948 37300
rect 77320 36800 77720 37300
rect 81092 36800 81492 37300
rect 84864 36800 85264 37300
rect 300 36400 97300 36800
rect 300 35800 13250 36200
rect 13550 35800 17022 36200
rect 17322 35800 20794 36200
rect 21094 35800 35882 36200
rect 36182 35800 47198 36200
rect 47498 35800 62286 36200
rect 62586 35800 66058 36200
rect 66358 35800 88690 36200
rect 88990 35800 92462 36200
rect 92762 35800 96234 36200
rect 96534 35800 97300 36200
rect 27310 34758 27550 34768
rect 23220 34748 24260 34758
rect 23450 34568 24260 34748
rect 23220 34368 24260 34568
rect 27310 34138 27320 34758
rect 27540 34368 28140 34758
rect 27540 34138 27550 34368
rect 27310 33938 27550 34138
rect 1880 32178 2280 33038
rect 5652 32178 6052 32678
rect 9424 32178 9824 32678
rect 24512 32178 24912 32678
rect 28284 32178 28684 32678
rect 32056 32178 32456 32678
rect 39600 32178 40000 32678
rect 43372 32178 43772 32678
rect 50916 32178 51316 32678
rect 54688 32178 55088 32678
rect 58460 32178 58860 32678
rect 69776 32178 70176 32678
rect 73548 32178 73948 32678
rect 77320 32178 77720 32678
rect 81092 32178 81492 32678
rect 84864 32178 85264 32678
rect 300 31778 97300 32178
rect 300 31178 13250 31578
rect 13550 31178 17022 31578
rect 17322 31178 20794 31578
rect 21094 31178 35882 31578
rect 36182 31178 47198 31578
rect 47498 31178 62286 31578
rect 62586 31178 66058 31578
rect 66358 31178 88690 31578
rect 88990 31178 92462 31578
rect 92762 31178 96234 31578
rect 96534 31178 97300 31578
rect 27310 30136 27550 30146
rect 23220 30126 24260 30136
rect 23450 29946 24260 30126
rect 23220 29746 24260 29946
rect 27310 29516 27320 30136
rect 27540 29746 28140 30136
rect 27540 29516 27550 29746
rect 27310 29316 27550 29516
rect 1880 27556 2280 28416
rect 5652 27556 6052 28056
rect 9424 27556 9824 28056
rect 24512 27556 24912 28056
rect 28284 27556 28684 28056
rect 32056 27556 32456 28056
rect 39600 27556 40000 28056
rect 43372 27556 43772 28056
rect 50916 27556 51316 28056
rect 54688 27556 55088 28056
rect 58460 27556 58860 28056
rect 69776 27556 70176 28056
rect 73548 27556 73948 28056
rect 77320 27556 77720 28056
rect 81092 27556 81492 28056
rect 84864 27556 85264 28056
rect 300 27156 97300 27556
rect 300 26556 13250 26956
rect 13550 26556 17022 26956
rect 17322 26556 20794 26956
rect 21094 26556 35882 26956
rect 36182 26556 47198 26956
rect 47498 26556 62286 26956
rect 62586 26556 66058 26956
rect 66358 26556 88690 26956
rect 88990 26556 92462 26956
rect 92762 26556 96234 26956
rect 96534 26556 97300 26956
rect 27310 25514 27550 25524
rect 23220 25504 24260 25514
rect 23450 25324 24260 25504
rect 23220 25124 24260 25324
rect 27310 24894 27320 25514
rect 27540 25124 28140 25514
rect 27540 24894 27550 25124
rect 27310 24694 27550 24894
rect 1880 22934 2280 23794
rect 5652 22934 6052 23434
rect 9424 22934 9824 23434
rect 24512 22934 24912 23434
rect 28284 22934 28684 23434
rect 32056 22934 32456 23434
rect 39600 22934 40000 23434
rect 54688 22934 55088 23434
rect 58460 22934 58860 23434
rect 73548 22934 73948 23434
rect 77320 22934 77720 23434
rect 81092 22934 81492 23434
rect 84864 22934 85264 23434
rect 300 22534 97300 22934
rect 300 21934 13250 22334
rect 13550 21934 17022 22334
rect 17322 21934 20794 22334
rect 21094 21934 35882 22334
rect 36182 21934 47198 22334
rect 47498 21934 62286 22334
rect 62586 21934 66058 22334
rect 66358 21934 88690 22334
rect 88990 21934 92462 22334
rect 92762 21934 96234 22334
rect 96534 21934 97300 22334
rect 39460 21340 43426 21740
rect 43726 21340 50970 21740
rect 51270 21340 69830 21740
rect 70130 21340 71780 21740
rect 27310 20892 27550 20902
rect 23220 20882 24260 20892
rect 23450 20702 24260 20882
rect 23220 20502 24260 20702
rect 27310 20272 27320 20892
rect 27540 20502 28140 20892
rect 27540 20272 27550 20502
rect 27310 20072 27550 20272
rect 1880 18312 2280 19172
rect 5652 18312 6052 18812
rect 9424 18312 9824 18812
rect 24512 18312 24912 18812
rect 28284 18312 28684 18812
rect 32056 18312 32456 18812
rect 39600 18312 40000 18812
rect 54688 18312 55088 18812
rect 58460 18312 58860 18812
rect 73548 18312 73948 18812
rect 77320 18312 77720 18812
rect 81092 18312 81492 18812
rect 84864 18312 85264 18812
rect 300 17912 97300 18312
rect 300 17312 13250 17712
rect 13550 17312 17022 17712
rect 17322 17312 20794 17712
rect 21094 17312 35882 17712
rect 36182 17312 47198 17712
rect 47498 17312 62286 17712
rect 62586 17312 66058 17712
rect 66358 17312 88690 17712
rect 88990 17312 92462 17712
rect 92762 17312 96234 17712
rect 96534 17312 97300 17712
rect 39460 16718 43426 17118
rect 43726 16718 50970 17118
rect 51270 16718 69830 17118
rect 70130 16718 71780 17118
rect 27310 16270 27550 16280
rect 23220 16260 24490 16270
rect 23450 16080 24490 16260
rect 23220 15880 24490 16080
rect 27310 15650 27320 16270
rect 27540 15880 28140 16270
rect 27540 15650 27550 15880
rect 27310 15450 27550 15650
rect 1880 13690 2280 14550
rect 5652 13690 6052 14190
rect 9424 13690 9824 14190
rect 24512 13690 24912 14190
rect 28284 13690 28684 14190
rect 32056 13690 32456 14190
rect 39600 13690 40000 14190
rect 54688 13690 55088 14190
rect 58460 13690 58860 14190
rect 73548 13690 73948 14190
rect 77320 13690 77720 14190
rect 81092 13690 81492 14190
rect 84864 13690 85264 14190
rect 300 13290 97300 13690
rect 300 12690 13250 13090
rect 13550 12690 17022 13090
rect 17322 12690 20794 13090
rect 21094 12690 35882 13090
rect 36182 12690 47198 13090
rect 47498 12690 62286 13090
rect 62586 12690 66058 13090
rect 66358 12690 88690 13090
rect 88990 12690 92462 13090
rect 92762 12690 96234 13090
rect 96534 12690 97300 13090
rect 39460 12096 43426 12496
rect 43726 12096 50970 12496
rect 51270 12096 69830 12496
rect 70130 12096 71780 12496
rect 3110 9330 3380 9950
rect 4020 9330 4290 9950
rect 3110 9120 4290 9330
rect 18190 9330 18460 9550
rect 19110 9330 19380 9550
rect 18190 9120 19380 9330
rect 6960 8330 7620 8340
rect 3380 8250 3860 8260
rect 3380 7710 3390 8250
rect 3850 7900 3860 8250
rect 6960 7970 6970 8330
rect 7610 8180 7620 8330
rect 15740 8330 16400 8340
rect 15740 8190 15750 8330
rect 7610 7980 9890 8180
rect 7610 7970 7620 7980
rect 6960 7960 7620 7970
rect 3850 7890 9520 7900
rect 3850 7710 9260 7890
rect 3380 7700 9260 7710
rect 9250 7580 9260 7700
rect 9510 7580 9520 7890
rect 9250 7570 9520 7580
rect 9620 7890 9890 7980
rect 9620 7580 9630 7890
rect 9880 7580 9890 7890
rect 12950 7990 15750 8190
rect 12950 7900 13220 7990
rect 15740 7970 15750 7990
rect 16390 7970 16400 8330
rect 15740 7960 16400 7970
rect 19510 8320 19990 8330
rect 12950 7590 12960 7900
rect 13210 7590 13220 7900
rect 12950 7580 13220 7590
rect 13320 7900 13590 7910
rect 19510 7900 19520 8320
rect 13320 7590 13330 7900
rect 13580 7780 19520 7900
rect 19980 7780 19990 8320
rect 13580 7700 19990 7780
rect 13580 7590 13590 7700
rect 13320 7580 13590 7590
rect 9620 7570 9890 7580
rect 8200 7190 8920 7200
rect 8200 6710 8220 7190
rect 8900 6710 8920 7190
rect 8200 6700 8920 6710
rect 12000 7190 12700 7200
rect 12000 6710 12010 7190
rect 12690 6710 12700 7190
rect 47960 6860 47980 7050
rect 12000 6700 12700 6710
rect 43310 6670 47980 6860
rect 48350 6670 48370 7050
rect 43310 6660 48370 6670
rect 43310 6460 43530 6660
rect 52330 6610 52730 6620
rect 39440 6450 43530 6460
rect 39440 6270 39450 6450
rect 41650 6270 43530 6450
rect 39440 6260 43530 6270
rect 44790 6410 45190 6460
rect 44790 6030 44800 6410
rect 45180 6030 45190 6410
rect 47840 6450 50060 6460
rect 47840 6270 47850 6450
rect 50050 6270 50060 6450
rect 52330 6420 52340 6610
rect 47840 6260 50060 6270
rect 50720 6410 52340 6420
rect 50720 6230 50730 6410
rect 51280 6230 52340 6410
rect 52720 6230 52730 6610
rect 50720 6220 52730 6230
rect 44790 6020 45190 6030
rect 37950 5790 45930 5800
rect 9100 5440 9260 5450
rect 9100 5140 9110 5440
rect 9250 5350 9260 5440
rect 9530 5440 9610 5450
rect 9530 5350 9540 5440
rect 9250 5150 9540 5350
rect 9250 5140 9260 5150
rect 9100 5130 9260 5140
rect 9530 5140 9540 5150
rect 9600 5350 9610 5440
rect 9880 5440 10040 5450
rect 9880 5350 9890 5440
rect 9600 5150 9890 5350
rect 9600 5140 9610 5150
rect 9530 5130 9610 5140
rect 9880 5140 9890 5150
rect 10030 5350 10040 5440
rect 12800 5440 12960 5450
rect 10240 5350 10650 5360
rect 10030 5150 10250 5350
rect 10030 5140 10040 5150
rect 9880 5130 10040 5140
rect 9100 4800 9260 4810
rect 9100 4500 9110 4800
rect 9250 4790 9260 4800
rect 9530 4800 9610 4810
rect 9530 4790 9540 4800
rect 9250 4590 9540 4790
rect 9250 4500 9260 4590
rect 9100 4490 9260 4500
rect 9530 4500 9540 4590
rect 9600 4790 9610 4800
rect 9880 4800 10040 4810
rect 9880 4790 9890 4800
rect 9600 4590 9890 4790
rect 9600 4500 9610 4590
rect 9530 4490 9610 4500
rect 9880 4500 9890 4590
rect 10030 4790 10040 4800
rect 10240 4790 10250 5150
rect 10030 4590 10250 4790
rect 10640 4590 10650 5350
rect 12800 5140 12810 5440
rect 12950 5350 12960 5440
rect 13230 5440 13310 5450
rect 13230 5350 13240 5440
rect 12950 5150 13240 5350
rect 12950 5140 12960 5150
rect 12800 5130 12960 5140
rect 13230 5140 13240 5150
rect 13300 5350 13310 5440
rect 13590 5440 13750 5450
rect 13590 5350 13600 5440
rect 13300 5150 13600 5350
rect 13300 5140 13310 5150
rect 13230 5130 13310 5140
rect 13590 5140 13600 5150
rect 13740 5350 13750 5440
rect 37950 5410 37960 5790
rect 38270 5410 39240 5790
rect 39410 5410 39690 5790
rect 39750 5410 40010 5790
rect 40070 5410 40330 5790
rect 40390 5410 40640 5790
rect 40700 5410 40960 5790
rect 41020 5410 41270 5790
rect 41330 5410 41590 5790
rect 41650 5410 41940 5790
rect 42110 5410 45540 5790
rect 45920 5410 45930 5790
rect 37950 5400 45930 5410
rect 47630 5790 50530 5800
rect 47630 5410 47640 5790
rect 47810 5410 48090 5790
rect 48150 5410 48410 5790
rect 48470 5410 48730 5790
rect 48790 5410 49040 5790
rect 49100 5410 49360 5790
rect 49420 5410 49670 5790
rect 49730 5410 49990 5790
rect 50050 5410 50340 5790
rect 50510 5410 50530 5790
rect 47630 5400 50530 5410
rect 14010 5350 14420 5360
rect 13740 5150 14020 5350
rect 13740 5140 13750 5150
rect 13590 5130 13750 5140
rect 10030 4500 10040 4590
rect 10240 4580 10650 4590
rect 12800 4800 12960 4810
rect 9880 4490 10040 4500
rect 12800 4500 12810 4800
rect 12950 4790 12960 4800
rect 13230 4800 13310 4810
rect 13230 4790 13240 4800
rect 12950 4590 13240 4790
rect 12950 4500 12960 4590
rect 12800 4490 12960 4500
rect 13230 4500 13240 4590
rect 13300 4790 13310 4800
rect 13590 4800 13750 4810
rect 13590 4790 13600 4800
rect 13300 4590 13600 4790
rect 13300 4500 13310 4590
rect 13230 4490 13310 4500
rect 13590 4500 13600 4590
rect 13740 4790 13750 4800
rect 14010 4790 14020 5150
rect 13740 4590 14020 4790
rect 14410 4590 14420 5350
rect 44190 5190 44590 5200
rect 38620 5040 38870 5050
rect 13740 4500 13750 4590
rect 14010 4580 14420 4590
rect 13590 4490 13750 4500
rect 9370 4480 9450 4490
rect 6460 4310 8860 4320
rect 6460 4130 6480 4310
rect 6860 4130 8570 4310
rect 8850 4130 8860 4310
rect 6460 4120 8860 4130
rect 9370 4000 9380 4480
rect 2700 3990 9380 4000
rect 2700 3810 2710 3990
rect 3090 3880 9380 3990
rect 9440 3880 9450 4480
rect 3090 3810 9450 3880
rect 2700 3800 9450 3810
rect 13390 4480 13470 4490
rect 13390 3810 13400 4480
rect 13460 4000 13470 4480
rect 38620 4420 38630 5040
rect 38860 4420 38870 5040
rect 39440 4940 41820 4950
rect 39440 4760 39450 4940
rect 41810 4760 41820 4940
rect 44190 4810 44200 5190
rect 44580 4810 44590 5190
rect 51730 5190 52130 5200
rect 51730 5000 51740 5190
rect 50710 4990 51740 5000
rect 44190 4800 44590 4810
rect 47840 4940 50220 4950
rect 39440 4750 40430 4760
rect 40420 4560 40430 4750
rect 40810 4750 41820 4760
rect 47840 4760 47850 4940
rect 50210 4760 50220 4940
rect 50710 4810 50720 4990
rect 51270 4810 51740 4990
rect 52120 4810 52130 5190
rect 50710 4800 52130 4810
rect 47840 4750 50220 4760
rect 40810 4560 40820 4750
rect 40420 4550 40820 4560
rect 38620 4410 38870 4420
rect 13960 4310 17790 4320
rect 13960 4130 13970 4310
rect 14250 4130 17790 4310
rect 13960 4120 17790 4130
rect 18180 4120 18200 4320
rect 43860 4280 47800 4290
rect 37410 4250 40960 4260
rect 13460 3810 21570 4000
rect 13390 3800 21570 3810
rect 21950 3800 21960 4000
rect 37410 3870 37420 4250
rect 37790 3870 40770 4250
rect 40950 3870 40960 4250
rect 43860 4100 43870 4280
rect 44580 4100 47490 4280
rect 47790 4100 47800 4280
rect 43860 4090 47800 4100
rect 51920 4230 52310 4240
rect 51920 4020 51930 4230
rect 37410 3860 40960 3870
rect 44380 4010 51930 4020
rect 44380 3830 44390 4010
rect 45100 3830 51930 4010
rect 52300 3830 52310 4230
rect 44380 3820 52310 3830
rect 44890 3740 56660 3750
rect 36640 3720 39930 3730
rect 36640 3340 36650 3720
rect 37040 3340 39740 3720
rect 39920 3340 39930 3720
rect 44890 3560 44900 3740
rect 45610 3560 56280 3740
rect 44890 3550 56280 3560
rect 36640 3330 39930 3340
rect 56270 3340 56280 3550
rect 56650 3340 56660 3740
rect 56270 3330 56660 3340
rect 33640 3230 40450 3240
rect 33640 2850 33650 3230
rect 34020 2850 40260 3230
rect 40440 2850 40450 3230
rect 33640 2840 40450 2850
rect 38220 2690 46060 2700
rect 38220 2310 38230 2690
rect 38610 2310 38770 2690
rect 38830 2310 39030 2690
rect 39090 2310 39540 2690
rect 39600 2310 40060 2690
rect 40120 2310 40580 2690
rect 40640 2310 41090 2690
rect 41150 2310 41610 2690
rect 41670 2310 42120 2690
rect 42180 2310 42640 2690
rect 42700 2310 43160 2690
rect 43220 2310 43670 2690
rect 43730 2310 44190 2690
rect 44250 2310 44700 2690
rect 44760 2310 45220 2690
rect 45280 2310 45740 2690
rect 45800 2310 45990 2690
rect 46050 2310 46060 2690
rect 38220 2300 46060 2310
rect 32640 2230 45750 2240
rect 32640 2110 39100 2230
rect 39240 2110 39400 2230
rect 39750 2110 39910 2230
rect 40260 2110 40430 2230
rect 40780 2110 40940 2230
rect 41290 2110 41460 2230
rect 41810 2110 41980 2230
rect 42330 2110 42490 2230
rect 42840 2110 43010 2230
rect 43360 2110 43520 2230
rect 43870 2110 44040 2230
rect 44390 2110 44560 2230
rect 44910 2110 45070 2230
rect 45420 2110 45590 2230
rect 45730 2110 45750 2230
rect 32640 2100 45750 2110
rect 32870 1990 39420 2000
rect 32870 1610 32880 1990
rect 33270 1610 39230 1990
rect 39410 1610 39420 1990
rect 32870 1600 39420 1610
rect 38220 1470 46060 1480
rect 38220 1090 38230 1470
rect 38610 1090 38770 1470
rect 38830 1090 39030 1470
rect 39090 1090 39540 1470
rect 39600 1090 40060 1470
rect 40120 1090 40580 1470
rect 40640 1090 41090 1470
rect 41150 1090 41610 1470
rect 41670 1090 42120 1470
rect 42180 1090 42640 1470
rect 42700 1090 43160 1470
rect 43220 1090 43670 1470
rect 43730 1090 44190 1470
rect 44250 1090 44700 1470
rect 44760 1090 45220 1470
rect 45280 1090 45740 1470
rect 45800 1090 45990 1470
rect 46050 1090 46060 1470
rect 38220 1080 46060 1090
rect 33640 960 39930 970
rect 33640 580 33650 960
rect 34010 580 39740 960
rect 39920 580 39930 960
rect 33640 570 39930 580
<< via3 >>
rect 2710 38990 3094 39374
rect 6482 38990 6866 39374
rect 10254 38990 10638 39374
rect 14026 38990 14410 39374
rect 17798 38990 18182 39374
rect 21570 38990 21954 39374
rect 23220 39190 23450 39370
rect 25342 38990 25726 39374
rect 27320 38760 27540 39380
rect 29114 38990 29498 39374
rect 32886 38990 33270 39374
rect 36658 38990 37042 39374
rect 40430 38990 40814 39374
rect 44202 38990 44586 39374
rect 47974 38990 48358 39374
rect 51746 38990 52130 39374
rect 55518 38990 55902 39374
rect 59290 38990 59674 39374
rect 63062 38990 63446 39374
rect 66834 38990 67218 39374
rect 70606 38990 70990 39374
rect 74378 38990 74762 39374
rect 78150 38990 78534 39374
rect 81922 38990 82306 39374
rect 85694 38990 86078 39374
rect 89466 38990 89850 39374
rect 93238 38990 93622 39374
rect 97010 38990 97394 39374
rect 13250 35800 13550 36200
rect 17022 35800 17322 36200
rect 20794 35800 21094 36200
rect 35882 35800 36182 36200
rect 47198 35800 47498 36200
rect 62286 35800 62586 36200
rect 66058 35800 66358 36200
rect 88690 35800 88990 36200
rect 92462 35800 92762 36200
rect 96234 35800 96534 36200
rect 2710 34368 3094 34752
rect 6482 34368 6866 34752
rect 10254 34368 10638 34752
rect 14026 34368 14410 34752
rect 17798 34368 18182 34752
rect 21570 34368 21954 34752
rect 23220 34568 23450 34748
rect 25342 34368 25726 34752
rect 27320 34138 27540 34758
rect 29114 34368 29498 34752
rect 32886 34368 33270 34752
rect 36658 34368 37042 34752
rect 40430 34368 40814 34752
rect 44202 34368 44586 34752
rect 47974 34368 48358 34752
rect 51746 34368 52130 34752
rect 55518 34368 55902 34752
rect 59290 34368 59674 34752
rect 63062 34368 63446 34752
rect 66834 34368 67218 34752
rect 70606 34368 70990 34752
rect 74378 34368 74762 34752
rect 78150 34368 78534 34752
rect 81922 34368 82306 34752
rect 85694 34368 86078 34752
rect 89466 34368 89850 34752
rect 93238 34368 93622 34752
rect 97010 34368 97394 34752
rect 13250 31178 13550 31578
rect 17022 31178 17322 31578
rect 20794 31178 21094 31578
rect 35882 31178 36182 31578
rect 47198 31178 47498 31578
rect 62286 31178 62586 31578
rect 66058 31178 66358 31578
rect 88690 31178 88990 31578
rect 92462 31178 92762 31578
rect 96234 31178 96534 31578
rect 2710 29746 3094 30130
rect 6482 29746 6866 30130
rect 10254 29746 10638 30130
rect 14026 29746 14410 30130
rect 17798 29746 18182 30130
rect 21570 29746 21954 30130
rect 23220 29946 23450 30126
rect 25342 29746 25726 30130
rect 27320 29516 27540 30136
rect 29114 29746 29498 30130
rect 32886 29746 33270 30130
rect 36658 29746 37042 30130
rect 40430 29746 40814 30130
rect 44202 29746 44586 30130
rect 47974 29746 48358 30130
rect 51746 29746 52130 30130
rect 55518 29746 55902 30130
rect 59290 29746 59674 30130
rect 63062 29746 63446 30130
rect 66834 29746 67218 30130
rect 70606 29746 70990 30130
rect 74378 29746 74762 30130
rect 78150 29746 78534 30130
rect 81922 29746 82306 30130
rect 85694 29746 86078 30130
rect 89466 29746 89850 30130
rect 93238 29746 93622 30130
rect 97010 29746 97394 30130
rect 13250 26556 13550 26956
rect 17022 26556 17322 26956
rect 20794 26556 21094 26956
rect 35882 26556 36182 26956
rect 47198 26556 47498 26956
rect 62286 26556 62586 26956
rect 66058 26556 66358 26956
rect 88690 26556 88990 26956
rect 92462 26556 92762 26956
rect 96234 26556 96534 26956
rect 2710 25124 3094 25508
rect 6482 25124 6866 25508
rect 10254 25124 10638 25508
rect 14026 25124 14410 25508
rect 17798 25124 18182 25508
rect 21570 25124 21954 25508
rect 23220 25324 23450 25504
rect 25342 25124 25726 25508
rect 27320 24894 27540 25514
rect 29114 25124 29498 25508
rect 32886 25124 33270 25508
rect 36658 25124 37042 25508
rect 40430 25124 40814 25508
rect 44802 25124 45186 25508
rect 47974 25124 48358 25508
rect 52346 25124 52730 25508
rect 55518 25124 55902 25508
rect 59290 25124 59674 25508
rect 63062 25124 63446 25508
rect 66834 25124 67218 25508
rect 71206 25124 71590 25508
rect 74378 25124 74762 25508
rect 78150 25124 78534 25508
rect 81922 25124 82306 25508
rect 85694 25124 86078 25508
rect 89466 25124 89850 25508
rect 93238 25124 93622 25508
rect 97010 25124 97394 25508
rect 13250 21934 13550 22334
rect 17022 21934 17322 22334
rect 20794 21934 21094 22334
rect 35882 21934 36182 22334
rect 47198 21934 47498 22334
rect 62286 21934 62586 22334
rect 66058 21934 66358 22334
rect 88690 21934 88990 22334
rect 92462 21934 92762 22334
rect 96234 21934 96534 22334
rect 43426 21340 43726 21740
rect 50970 21340 51270 21740
rect 69830 21340 70130 21740
rect 2710 20502 3094 20886
rect 6482 20502 6866 20886
rect 10254 20502 10638 20886
rect 14026 20502 14410 20886
rect 17798 20502 18182 20886
rect 21570 20502 21954 20886
rect 23220 20702 23450 20882
rect 25342 20502 25726 20886
rect 27320 20272 27540 20892
rect 29114 20502 29498 20886
rect 32886 20502 33270 20886
rect 36658 20502 37042 20886
rect 40430 20502 40814 20886
rect 44802 20502 45186 20886
rect 47974 20502 48358 20886
rect 52346 20502 52730 20886
rect 55518 20502 55902 20886
rect 59290 20502 59674 20886
rect 63062 20502 63446 20886
rect 66834 20502 67218 20886
rect 71206 20502 71590 20886
rect 74378 20502 74762 20886
rect 78150 20502 78534 20886
rect 81922 20502 82306 20886
rect 85694 20502 86078 20886
rect 89466 20502 89850 20886
rect 93238 20502 93622 20886
rect 97010 20502 97394 20886
rect 13250 17312 13550 17712
rect 17022 17312 17322 17712
rect 20794 17312 21094 17712
rect 35882 17312 36182 17712
rect 47198 17312 47498 17712
rect 62286 17312 62586 17712
rect 66058 17312 66358 17712
rect 88690 17312 88990 17712
rect 92462 17312 92762 17712
rect 96234 17312 96534 17712
rect 43426 16718 43726 17118
rect 50970 16718 51270 17118
rect 69830 16718 70130 17118
rect 2710 15880 3094 16264
rect 6482 15880 6866 16264
rect 10254 15880 10638 16264
rect 14026 15880 14410 16264
rect 17798 15880 18182 16264
rect 21570 15880 21954 16264
rect 23220 16080 23450 16260
rect 25342 15880 25726 16264
rect 27320 15650 27540 16270
rect 29114 15880 29498 16264
rect 32886 15880 33270 16264
rect 36658 15880 37042 16264
rect 40430 15880 40814 16264
rect 44802 15880 45186 16264
rect 47974 15880 48358 16264
rect 52346 15880 52730 16264
rect 55518 15880 55902 16264
rect 59290 15880 59674 16264
rect 63062 15880 63446 16264
rect 66834 15880 67218 16264
rect 71206 15880 71590 16264
rect 74378 15880 74762 16264
rect 78150 15880 78534 16264
rect 81922 15880 82306 16264
rect 85694 15880 86078 16264
rect 89466 15880 89850 16264
rect 93238 15880 93622 16264
rect 97010 15880 97394 16264
rect 13250 12690 13550 13090
rect 17022 12690 17322 13090
rect 20794 12690 21094 13090
rect 35882 12690 36182 13090
rect 47198 12690 47498 13090
rect 62286 12690 62586 13090
rect 66058 12690 66358 13090
rect 88690 12690 88990 13090
rect 92462 12690 92762 13090
rect 96234 12690 96534 13090
rect 43426 12096 43726 12496
rect 50970 12096 51270 12496
rect 69830 12096 70130 12496
rect 10250 11260 10640 11650
rect 14020 11260 14410 11650
rect 2710 9560 3090 9940
rect 8130 9550 8370 9940
rect 11900 9550 12140 9940
rect 32880 9550 33270 9940
rect 33650 9430 34020 9930
rect 36650 9550 37040 9940
rect 37420 9430 37790 9930
rect 8460 6710 8680 7180
rect 12230 6720 12450 7180
rect 47980 6670 48350 7050
rect 44800 6030 45180 6410
rect 52340 6230 52720 6610
rect 10250 4590 10640 5350
rect 14020 4590 14410 5350
rect 32880 4930 33270 5320
rect 36650 4930 37040 5320
rect 6480 4130 6860 4310
rect 2710 3810 3090 3990
rect 38630 4420 38860 5040
rect 40430 4760 40810 4940
rect 44200 4810 44580 5190
rect 40430 4560 40810 4760
rect 51740 4810 52120 5190
rect 17790 4120 18180 4320
rect 21570 3800 21950 4000
rect 37420 3870 37790 4250
rect 36650 3340 37040 3720
rect 33650 2850 34020 3230
rect 38230 2310 38610 2690
rect 32880 1610 33270 1990
rect 38230 1090 38610 1470
<< metal4 >>
rect 3006 44952 3066 45152
rect 3558 44952 3618 45152
rect 4110 44952 4170 45152
rect 4662 44952 4722 45152
rect 5214 44952 5274 45152
rect 5766 44952 5826 45152
rect 6318 44952 6378 45152
rect 6870 44952 6930 45152
rect 7422 44952 7482 45152
rect 7974 44952 8034 45152
rect 8526 44952 8586 45152
rect 9078 44952 9138 45152
rect 9630 44952 9690 45152
rect 10182 44952 10242 45152
rect 10734 44952 10794 45152
rect 11286 44952 11346 45152
rect 11838 44952 11898 45152
rect 12390 44952 12450 45152
rect 12942 44952 13002 45152
rect 13494 44952 13554 45152
rect 14046 44952 14106 45152
rect 14598 44952 14658 45152
rect 15150 44952 15210 45152
rect 15702 44952 15762 45152
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 44952 20730 45152
rect 21222 44952 21282 45152
rect 21774 44952 21834 45152
rect 22326 44952 22386 45152
rect 22878 44952 22938 45152
rect 23430 44952 23490 45152
rect 23982 44952 24042 45152
rect 24534 44952 24594 45152
rect 25086 44952 25146 45152
rect 25638 44952 25698 45152
rect 26190 44952 26250 45152
rect 2700 39374 3100 39600
rect 2700 38990 2710 39374
rect 3094 38990 3100 39374
rect 2700 34752 3100 38990
rect 2700 34368 2710 34752
rect 3094 34368 3100 34752
rect 2700 30130 3100 34368
rect 2700 29746 2710 30130
rect 3094 29746 3100 30130
rect 2700 25508 3100 29746
rect 2700 25124 2710 25508
rect 3094 25124 3100 25508
rect 2700 20886 3100 25124
rect 2700 20502 2710 20886
rect 3094 20502 3100 20886
rect 2700 16264 3100 20502
rect 2700 15880 2710 16264
rect 3094 15880 3100 16264
rect 2700 9940 3100 15880
rect 2700 9560 2710 9940
rect 3090 9560 3100 9940
rect 2700 3990 3100 9560
rect 2700 3810 2710 3990
rect 3090 3810 3100 3990
rect 2700 2980 3100 3810
rect 6472 39374 6872 39600
rect 6472 38990 6482 39374
rect 6866 38990 6872 39374
rect 6472 34752 6872 38990
rect 6472 34368 6482 34752
rect 6866 34368 6872 34752
rect 6472 30130 6872 34368
rect 6472 29746 6482 30130
rect 6866 29746 6872 30130
rect 6472 25508 6872 29746
rect 6472 25124 6482 25508
rect 6866 25124 6872 25508
rect 6472 20886 6872 25124
rect 6472 20502 6482 20886
rect 6866 20502 6872 20886
rect 6472 16264 6872 20502
rect 6472 15880 6482 16264
rect 6866 15880 6872 16264
rect 6472 4310 6872 15880
rect 10244 39374 10644 39600
rect 10244 38990 10254 39374
rect 10638 38990 10644 39374
rect 10244 34752 10644 38990
rect 14016 39374 14416 39600
rect 14016 38990 14026 39374
rect 14410 38990 14416 39374
rect 13300 36210 13500 38090
rect 13240 36200 13560 36210
rect 13240 35800 13250 36200
rect 13550 35800 13560 36200
rect 13240 35790 13560 35800
rect 10244 34368 10254 34752
rect 10638 34368 10644 34752
rect 10244 30130 10644 34368
rect 14016 34752 14416 38990
rect 17788 39374 18188 39600
rect 17788 38990 17798 39374
rect 18182 38990 18188 39374
rect 17072 36210 17272 38090
rect 17012 36200 17332 36210
rect 17012 35800 17022 36200
rect 17322 35800 17332 36200
rect 17012 35790 17332 35800
rect 14016 34368 14026 34752
rect 14410 34368 14416 34752
rect 13300 31588 13500 33468
rect 13240 31578 13560 31588
rect 13240 31178 13250 31578
rect 13550 31178 13560 31578
rect 13240 31168 13560 31178
rect 10244 29746 10254 30130
rect 10638 29746 10644 30130
rect 10244 25508 10644 29746
rect 14016 30130 14416 34368
rect 17788 34752 18188 38990
rect 21560 39374 21960 39600
rect 21560 38990 21570 39374
rect 21954 38990 21960 39374
rect 25332 39374 25732 39600
rect 20844 36210 21044 38090
rect 20784 36200 21104 36210
rect 20784 35800 20794 36200
rect 21094 35800 21104 36200
rect 20784 35790 21104 35800
rect 17788 34368 17798 34752
rect 18182 34368 18188 34752
rect 17072 31588 17272 33468
rect 17012 31578 17332 31588
rect 17012 31178 17022 31578
rect 17322 31178 17332 31578
rect 17012 31168 17332 31178
rect 14016 29746 14026 30130
rect 14410 29746 14416 30130
rect 13300 26966 13500 28846
rect 13240 26956 13560 26966
rect 13240 26556 13250 26956
rect 13550 26556 13560 26956
rect 13240 26546 13560 26556
rect 10244 25124 10254 25508
rect 10638 25124 10644 25508
rect 10244 20886 10644 25124
rect 14016 25508 14416 29746
rect 17788 30130 18188 34368
rect 21560 34752 21960 38990
rect 21560 34368 21570 34752
rect 21954 34368 21960 34752
rect 25332 38990 25342 39374
rect 25726 38990 25732 39374
rect 25332 34752 25732 38990
rect 29104 39374 29504 39600
rect 29104 38990 29114 39374
rect 29498 38990 29504 39374
rect 20844 31588 21044 33468
rect 20784 31578 21104 31588
rect 20784 31178 20794 31578
rect 21094 31178 21104 31578
rect 20784 31168 21104 31178
rect 17788 29746 17798 30130
rect 18182 29746 18188 30130
rect 17072 26966 17272 28846
rect 17012 26956 17332 26966
rect 17012 26556 17022 26956
rect 17322 26556 17332 26956
rect 17012 26546 17332 26556
rect 14016 25124 14026 25508
rect 14410 25124 14416 25508
rect 13300 22344 13500 24224
rect 13240 22334 13560 22344
rect 13240 21934 13250 22334
rect 13550 21934 13560 22334
rect 13240 21924 13560 21934
rect 10244 20502 10254 20886
rect 10638 20502 10644 20886
rect 10244 16264 10644 20502
rect 14016 20886 14416 25124
rect 17788 25508 18188 29746
rect 21560 30130 21960 34368
rect 21560 29746 21570 30130
rect 21954 29746 21960 30130
rect 25332 34368 25342 34752
rect 25726 34368 25732 34752
rect 25332 30130 25732 34368
rect 29104 34752 29504 38990
rect 29104 34368 29114 34752
rect 29498 34368 29504 34752
rect 20844 26966 21044 28846
rect 20784 26956 21104 26966
rect 20784 26556 20794 26956
rect 21094 26556 21104 26956
rect 20784 26546 21104 26556
rect 17788 25124 17798 25508
rect 18182 25124 18188 25508
rect 17072 22344 17272 24224
rect 17012 22334 17332 22344
rect 17012 21934 17022 22334
rect 17322 21934 17332 22334
rect 17012 21924 17332 21934
rect 14016 20502 14026 20886
rect 14410 20502 14416 20886
rect 13300 17722 13500 19602
rect 13240 17712 13560 17722
rect 13240 17312 13250 17712
rect 13550 17312 13560 17712
rect 13240 17302 13560 17312
rect 10244 15880 10254 16264
rect 10638 15880 10644 16264
rect 10244 11650 10644 15880
rect 14016 16264 14416 20502
rect 17788 20886 18188 25124
rect 21560 25508 21960 29746
rect 21560 25124 21570 25508
rect 21954 25124 21960 25508
rect 25332 29746 25342 30130
rect 25726 29746 25732 30130
rect 25332 25508 25732 29746
rect 29104 30130 29504 34368
rect 29104 29746 29114 30130
rect 29498 29746 29504 30130
rect 20844 22344 21044 24224
rect 20784 22334 21104 22344
rect 20784 21934 20794 22334
rect 21094 21934 21104 22334
rect 20784 21924 21104 21934
rect 17788 20502 17798 20886
rect 18182 20502 18188 20886
rect 17072 17722 17272 19602
rect 17012 17712 17332 17722
rect 17012 17312 17022 17712
rect 17322 17312 17332 17712
rect 17012 17302 17332 17312
rect 14016 15880 14026 16264
rect 14410 15880 14416 16264
rect 13300 13100 13500 14980
rect 13240 13090 13560 13100
rect 13240 12690 13250 13090
rect 13550 12690 13560 13090
rect 13240 12680 13560 12690
rect 10244 11260 10250 11650
rect 10640 11260 10644 11650
rect 8120 9940 8380 9960
rect 8120 9550 8130 9940
rect 8370 9550 8380 9940
rect 8120 9540 8380 9550
rect 6472 4130 6480 4310
rect 6860 4130 6872 4310
rect 6472 2980 6872 4130
rect 10244 5350 10644 11260
rect 14016 11650 14416 15880
rect 17788 16264 18188 20502
rect 21560 20886 21960 25124
rect 21560 20502 21570 20886
rect 21954 20502 21960 20886
rect 25332 25124 25342 25508
rect 25726 25124 25732 25508
rect 25332 20886 25732 25124
rect 29104 25508 29504 29746
rect 29104 25124 29114 25508
rect 29498 25124 29504 25508
rect 20844 17722 21044 19602
rect 20784 17712 21104 17722
rect 20784 17312 20794 17712
rect 21094 17312 21104 17712
rect 20784 17302 21104 17312
rect 17788 15880 17798 16264
rect 18182 15880 18188 16264
rect 17072 13100 17272 14980
rect 17012 13090 17332 13100
rect 17012 12690 17022 13090
rect 17322 12690 17332 13090
rect 17012 12680 17332 12690
rect 14016 11260 14020 11650
rect 14410 11260 14416 11650
rect 11890 9940 12150 9960
rect 11890 9550 11900 9940
rect 12140 9550 12150 9940
rect 11890 9540 12150 9550
rect 10244 4590 10250 5350
rect 10640 4590 10644 5350
rect 10244 2980 10644 4590
rect 14016 5350 14416 11260
rect 14016 4590 14020 5350
rect 14410 4590 14416 5350
rect 14016 2980 14416 4590
rect 17788 4320 18188 15880
rect 21560 16264 21960 20502
rect 21560 15880 21570 16264
rect 21954 15880 21960 16264
rect 25332 20502 25342 20886
rect 25726 20502 25732 20886
rect 25332 16264 25732 20502
rect 29104 20886 29504 25124
rect 29104 20502 29114 20886
rect 29498 20502 29504 20886
rect 20844 13100 21044 14980
rect 20784 13090 21104 13100
rect 20784 12690 20794 13090
rect 21094 12690 21104 13090
rect 20784 12680 21104 12690
rect 17788 4120 17790 4320
rect 18180 4120 18188 4320
rect 17788 2980 18188 4120
rect 21560 4000 21960 15880
rect 25332 15880 25342 16264
rect 25726 15880 25732 16264
rect 25332 15000 25732 15880
rect 29104 16264 29504 20502
rect 29104 15880 29114 16264
rect 29498 15880 29504 16264
rect 29104 15000 29504 15880
rect 32876 39374 33276 39600
rect 32876 38990 32886 39374
rect 33270 38990 33276 39374
rect 32876 34752 33276 38990
rect 36648 39374 37048 39600
rect 36648 38990 36658 39374
rect 37042 38990 37048 39374
rect 35932 36210 36132 38090
rect 35870 36200 36190 36210
rect 35870 35800 35882 36200
rect 36182 35800 36190 36200
rect 35870 35790 36190 35800
rect 32876 34368 32886 34752
rect 33270 34368 33276 34752
rect 32876 30130 33276 34368
rect 36648 34752 37048 38990
rect 36648 34368 36658 34752
rect 37042 34368 37048 34752
rect 35932 31588 36132 33468
rect 35870 31578 36190 31588
rect 35870 31178 35882 31578
rect 36182 31178 36190 31578
rect 35870 31168 36190 31178
rect 32876 29746 32886 30130
rect 33270 29746 33276 30130
rect 32876 25508 33276 29746
rect 36648 30130 37048 34368
rect 36648 29746 36658 30130
rect 37042 29746 37048 30130
rect 35932 26966 36132 28846
rect 35870 26956 36190 26966
rect 35870 26556 35882 26956
rect 36182 26556 36190 26956
rect 35870 26546 36190 26556
rect 32876 25124 32886 25508
rect 33270 25124 33276 25508
rect 32876 20886 33276 25124
rect 36648 25508 37048 29746
rect 36648 25124 36658 25508
rect 37042 25124 37048 25508
rect 35932 22344 36132 24224
rect 35870 22334 36190 22344
rect 35870 21934 35882 22334
rect 36182 21934 36190 22334
rect 35870 21924 36190 21934
rect 32876 20502 32886 20886
rect 33270 20502 33276 20886
rect 32876 16264 33276 20502
rect 36648 20886 37048 25124
rect 36648 20502 36658 20886
rect 37042 20502 37048 20886
rect 35932 17722 36132 19602
rect 35870 17712 36190 17722
rect 35870 17312 35882 17712
rect 36182 17312 36190 17712
rect 35870 17302 36190 17312
rect 32876 15880 32886 16264
rect 33270 15880 33276 16264
rect 32876 15000 33276 15880
rect 36648 16264 37048 20502
rect 36648 15880 36658 16264
rect 37042 15880 37048 16264
rect 36648 15000 37048 15880
rect 40420 39374 40820 39600
rect 40420 38990 40430 39374
rect 40814 38990 40820 39374
rect 40420 34752 40820 38990
rect 40420 34368 40430 34752
rect 40814 34368 40820 34752
rect 40420 30130 40820 34368
rect 40420 29746 40430 30130
rect 40814 29746 40820 30130
rect 40420 25508 40820 29746
rect 40420 25124 40430 25508
rect 40814 25124 40820 25508
rect 40420 20886 40820 25124
rect 44192 39374 44592 39600
rect 44192 38990 44202 39374
rect 44586 38990 44592 39374
rect 44192 34752 44592 38990
rect 44192 34368 44202 34752
rect 44586 34368 44592 34752
rect 44192 30130 44592 34368
rect 44192 29746 44202 30130
rect 44586 29746 44592 30130
rect 43476 21750 43676 24224
rect 43414 21740 43734 21750
rect 43414 21340 43426 21740
rect 43726 21340 43734 21740
rect 43414 21330 43734 21340
rect 40420 20502 40430 20886
rect 40814 20502 40820 20886
rect 40420 16264 40820 20502
rect 43476 17128 43676 19602
rect 43414 17118 43734 17128
rect 43414 16718 43426 17118
rect 43726 16718 43734 17118
rect 43414 16708 43734 16718
rect 40420 15880 40430 16264
rect 40814 15880 40820 16264
rect 21560 3800 21570 4000
rect 21950 3800 21960 4000
rect 21560 2980 21960 3800
rect 32870 9940 33280 15000
rect 35932 13100 36132 14980
rect 35870 13090 36190 13100
rect 35870 12690 35882 13090
rect 36182 12690 36190 13090
rect 35870 12680 36190 12690
rect 36640 9940 37050 15000
rect 32870 9550 32880 9940
rect 33270 9550 33280 9940
rect 32870 5320 33280 9550
rect 32870 4930 32880 5320
rect 33270 4930 33280 5320
rect 32870 1990 33280 4930
rect 33640 9930 34030 9940
rect 33640 9430 33650 9930
rect 34020 9430 34030 9930
rect 33640 3230 34030 9430
rect 33640 2850 33650 3230
rect 34020 2850 34030 3230
rect 33640 2840 34030 2850
rect 36640 9550 36650 9940
rect 37040 9550 37050 9940
rect 36640 5320 37050 9550
rect 36640 4930 36650 5320
rect 37040 4930 37050 5320
rect 36640 3720 37050 4930
rect 37410 9930 37800 9940
rect 37410 9430 37420 9930
rect 37790 9430 37800 9930
rect 37410 4250 37800 9430
rect 38620 5040 38870 5050
rect 38620 4420 38630 5040
rect 38860 4420 38870 5040
rect 40420 4940 40820 15880
rect 43476 12506 43676 14980
rect 43414 12496 43734 12506
rect 43414 12096 43426 12496
rect 43726 12096 43734 12496
rect 43414 12086 43734 12096
rect 44192 5200 44592 29746
rect 44792 25508 45192 39600
rect 47964 39374 48364 39600
rect 47964 38990 47974 39374
rect 48358 38990 48364 39374
rect 47248 36210 47448 38090
rect 47186 36200 47506 36210
rect 47186 35800 47198 36200
rect 47498 35800 47506 36200
rect 47186 35790 47506 35800
rect 47964 34752 48364 38990
rect 47964 34368 47974 34752
rect 48358 34368 48364 34752
rect 47248 31588 47448 33468
rect 47186 31578 47506 31588
rect 47186 31178 47198 31578
rect 47498 31178 47506 31578
rect 47186 31168 47506 31178
rect 47964 30130 48364 34368
rect 47964 29746 47974 30130
rect 48358 29746 48364 30130
rect 47248 26966 47448 28846
rect 47186 26956 47506 26966
rect 47186 26556 47198 26956
rect 47498 26556 47506 26956
rect 47186 26546 47506 26556
rect 44792 25124 44802 25508
rect 45186 25124 45192 25508
rect 44792 20886 45192 25124
rect 47964 25508 48364 29746
rect 47964 25124 47974 25508
rect 48358 25124 48364 25508
rect 47248 22344 47448 24224
rect 47186 22334 47506 22344
rect 47186 21934 47198 22334
rect 47498 21934 47506 22334
rect 47186 21924 47506 21934
rect 44792 20502 44802 20886
rect 45186 20502 45192 20886
rect 44792 16264 45192 20502
rect 47964 20886 48364 25124
rect 51736 39374 52136 39600
rect 51736 38990 51746 39374
rect 52130 38990 52136 39374
rect 51736 34752 52136 38990
rect 51736 34368 51746 34752
rect 52130 34368 52136 34752
rect 51736 30130 52136 34368
rect 51736 29746 51746 30130
rect 52130 29746 52136 30130
rect 51020 21750 51220 24224
rect 50958 21740 51278 21750
rect 50958 21340 50970 21740
rect 51270 21340 51278 21740
rect 50958 21330 51278 21340
rect 47964 20502 47974 20886
rect 48358 20502 48364 20886
rect 47248 17722 47448 19602
rect 47186 17712 47506 17722
rect 47186 17312 47198 17712
rect 47498 17312 47506 17712
rect 47186 17302 47506 17312
rect 44792 15880 44802 16264
rect 45186 15880 45192 16264
rect 44792 6420 45192 15880
rect 47964 16264 48364 20502
rect 51020 17128 51220 19602
rect 50958 17118 51278 17128
rect 50958 16718 50970 17118
rect 51270 16718 51278 17118
rect 50958 16708 51278 16718
rect 47964 15880 47974 16264
rect 48358 15880 48364 16264
rect 47248 13100 47448 14980
rect 47186 13090 47506 13100
rect 47186 12690 47198 13090
rect 47498 12690 47506 13090
rect 47186 12680 47506 12690
rect 47964 7050 48364 15880
rect 51020 12506 51220 14980
rect 50958 12496 51278 12506
rect 50958 12096 50970 12496
rect 51270 12096 51278 12496
rect 50958 12086 51278 12096
rect 47964 6670 47980 7050
rect 48350 6670 48364 7050
rect 47964 6660 48364 6670
rect 44790 6410 45192 6420
rect 44790 6030 44800 6410
rect 45180 6030 45192 6410
rect 44790 6020 45192 6030
rect 40420 4560 40430 4940
rect 40810 4560 40820 4940
rect 44190 5190 44592 5200
rect 44190 4810 44200 5190
rect 44580 4810 44592 5190
rect 44190 4800 44592 4810
rect 44792 4800 45192 6020
rect 51736 5200 52136 29746
rect 52336 25508 52736 39600
rect 52336 25124 52346 25508
rect 52730 25124 52736 25508
rect 52336 20886 52736 25124
rect 52336 20502 52346 20886
rect 52730 20502 52736 20886
rect 52336 16264 52736 20502
rect 52336 15880 52346 16264
rect 52730 15880 52736 16264
rect 52336 6620 52736 15880
rect 55508 39374 55908 39600
rect 55508 38990 55518 39374
rect 55902 38990 55908 39374
rect 55508 34752 55908 38990
rect 55508 34368 55518 34752
rect 55902 34368 55908 34752
rect 55508 30130 55908 34368
rect 55508 29746 55518 30130
rect 55902 29746 55908 30130
rect 55508 25508 55908 29746
rect 55508 25124 55518 25508
rect 55902 25124 55908 25508
rect 55508 20886 55908 25124
rect 55508 20502 55518 20886
rect 55902 20502 55908 20886
rect 55508 16264 55908 20502
rect 55508 15880 55518 16264
rect 55902 15880 55908 16264
rect 55508 15000 55908 15880
rect 59280 39374 59680 39600
rect 59280 38990 59290 39374
rect 59674 38990 59680 39374
rect 59280 34752 59680 38990
rect 63052 39374 63452 39600
rect 63052 38990 63062 39374
rect 63446 38990 63452 39374
rect 62336 36210 62536 38090
rect 62274 36200 62594 36210
rect 62274 35800 62286 36200
rect 62586 35800 62594 36200
rect 62274 35790 62594 35800
rect 59280 34368 59290 34752
rect 59674 34368 59680 34752
rect 59280 30130 59680 34368
rect 63052 34752 63452 38990
rect 66824 39374 67224 39600
rect 66824 38990 66834 39374
rect 67218 38990 67224 39374
rect 66108 36210 66308 38090
rect 66046 36200 66366 36210
rect 66046 35800 66058 36200
rect 66358 35800 66366 36200
rect 66046 35790 66366 35800
rect 63052 34368 63062 34752
rect 63446 34368 63452 34752
rect 62336 31588 62536 33468
rect 62274 31578 62594 31588
rect 62274 31178 62286 31578
rect 62586 31178 62594 31578
rect 62274 31168 62594 31178
rect 59280 29746 59290 30130
rect 59674 29746 59680 30130
rect 59280 25508 59680 29746
rect 63052 30130 63452 34368
rect 66824 34752 67224 38990
rect 66824 34368 66834 34752
rect 67218 34368 67224 34752
rect 66108 31588 66308 33468
rect 66046 31578 66366 31588
rect 66046 31178 66058 31578
rect 66358 31178 66366 31578
rect 66046 31168 66366 31178
rect 63052 29746 63062 30130
rect 63446 29746 63452 30130
rect 62336 26966 62536 28846
rect 62274 26956 62594 26966
rect 62274 26556 62286 26956
rect 62586 26556 62594 26956
rect 62274 26546 62594 26556
rect 59280 25124 59290 25508
rect 59674 25124 59680 25508
rect 59280 20886 59680 25124
rect 63052 25508 63452 29746
rect 66824 30130 67224 34368
rect 66824 29746 66834 30130
rect 67218 29746 67224 30130
rect 66108 26966 66308 28846
rect 66046 26956 66366 26966
rect 66046 26556 66058 26956
rect 66358 26556 66366 26956
rect 66046 26546 66366 26556
rect 63052 25124 63062 25508
rect 63446 25124 63452 25508
rect 62336 22344 62536 24224
rect 62274 22334 62594 22344
rect 62274 21934 62286 22334
rect 62586 21934 62594 22334
rect 62274 21924 62594 21934
rect 59280 20502 59290 20886
rect 59674 20502 59680 20886
rect 59280 16264 59680 20502
rect 63052 20886 63452 25124
rect 66824 25508 67224 29746
rect 66824 25124 66834 25508
rect 67218 25124 67224 25508
rect 66108 22344 66308 24224
rect 66046 22334 66366 22344
rect 66046 21934 66058 22334
rect 66358 21934 66366 22334
rect 66046 21924 66366 21934
rect 63052 20502 63062 20886
rect 63446 20502 63452 20886
rect 62336 17722 62536 19602
rect 62274 17712 62594 17722
rect 62274 17312 62286 17712
rect 62586 17312 62594 17712
rect 62274 17302 62594 17312
rect 59280 15880 59290 16264
rect 59674 15880 59680 16264
rect 59280 15000 59680 15880
rect 63052 16264 63452 20502
rect 66824 20886 67224 25124
rect 70596 39374 70996 39600
rect 70596 38990 70606 39374
rect 70990 38990 70996 39374
rect 70596 34752 70996 38990
rect 70596 34368 70606 34752
rect 70990 34368 70996 34752
rect 70596 30130 70996 34368
rect 70596 29746 70606 30130
rect 70990 29746 70996 30130
rect 69880 21750 70080 24224
rect 69818 21740 70138 21750
rect 69818 21340 69830 21740
rect 70130 21340 70138 21740
rect 69818 21330 70138 21340
rect 66824 20502 66834 20886
rect 67218 20502 67224 20886
rect 66108 17722 66308 19602
rect 66046 17712 66366 17722
rect 66046 17312 66058 17712
rect 66358 17312 66366 17712
rect 66046 17302 66366 17312
rect 63052 15880 63062 16264
rect 63446 15880 63452 16264
rect 63052 15000 63452 15880
rect 66824 16264 67224 20502
rect 69880 17128 70080 19602
rect 69818 17118 70138 17128
rect 69818 16718 69830 17118
rect 70130 16718 70138 17118
rect 69818 16708 70138 16718
rect 66824 15880 66834 16264
rect 67218 15880 67224 16264
rect 66824 15000 67224 15880
rect 70596 15000 70996 29746
rect 71196 25508 71596 39600
rect 71196 25124 71206 25508
rect 71590 25124 71596 25508
rect 71196 20886 71596 25124
rect 71196 20502 71206 20886
rect 71590 20502 71596 20886
rect 71196 16264 71596 20502
rect 71196 15880 71206 16264
rect 71590 15880 71596 16264
rect 71196 15000 71596 15880
rect 74368 39374 74768 39600
rect 74368 38990 74378 39374
rect 74762 38990 74768 39374
rect 74368 34752 74768 38990
rect 74368 34368 74378 34752
rect 74762 34368 74768 34752
rect 74368 30130 74768 34368
rect 74368 29746 74378 30130
rect 74762 29746 74768 30130
rect 74368 25508 74768 29746
rect 74368 25124 74378 25508
rect 74762 25124 74768 25508
rect 74368 20886 74768 25124
rect 74368 20502 74378 20886
rect 74762 20502 74768 20886
rect 74368 16264 74768 20502
rect 74368 15880 74378 16264
rect 74762 15880 74768 16264
rect 74368 15000 74768 15880
rect 78140 39374 78540 39600
rect 78140 38990 78150 39374
rect 78534 38990 78540 39374
rect 78140 34752 78540 38990
rect 78140 34368 78150 34752
rect 78534 34368 78540 34752
rect 78140 30130 78540 34368
rect 78140 29746 78150 30130
rect 78534 29746 78540 30130
rect 78140 25508 78540 29746
rect 78140 25124 78150 25508
rect 78534 25124 78540 25508
rect 78140 20886 78540 25124
rect 78140 20502 78150 20886
rect 78534 20502 78540 20886
rect 78140 16264 78540 20502
rect 78140 15880 78150 16264
rect 78534 15880 78540 16264
rect 78140 15000 78540 15880
rect 81912 39374 82312 39600
rect 81912 38990 81922 39374
rect 82306 38990 82312 39374
rect 81912 34752 82312 38990
rect 81912 34368 81922 34752
rect 82306 34368 82312 34752
rect 81912 30130 82312 34368
rect 81912 29746 81922 30130
rect 82306 29746 82312 30130
rect 81912 25508 82312 29746
rect 81912 25124 81922 25508
rect 82306 25124 82312 25508
rect 81912 20886 82312 25124
rect 81912 20502 81922 20886
rect 82306 20502 82312 20886
rect 81912 16264 82312 20502
rect 81912 15880 81922 16264
rect 82306 15880 82312 16264
rect 81912 15000 82312 15880
rect 85684 39374 86084 39600
rect 85684 38990 85694 39374
rect 86078 38990 86084 39374
rect 85684 34752 86084 38990
rect 89456 39374 89856 39600
rect 89456 38990 89466 39374
rect 89850 38990 89856 39374
rect 88740 36210 88940 38090
rect 88678 36200 88998 36210
rect 88678 35800 88690 36200
rect 88990 35800 88998 36200
rect 88678 35790 88998 35800
rect 85684 34368 85694 34752
rect 86078 34368 86084 34752
rect 85684 30130 86084 34368
rect 89456 34752 89856 38990
rect 93228 39374 93628 39600
rect 93228 38990 93238 39374
rect 93622 38990 93628 39374
rect 92512 36210 92712 38090
rect 92450 36200 92770 36210
rect 92450 35800 92462 36200
rect 92762 35800 92770 36200
rect 92450 35790 92770 35800
rect 89456 34368 89466 34752
rect 89850 34368 89856 34752
rect 88740 31588 88940 33468
rect 88678 31578 88998 31588
rect 88678 31178 88690 31578
rect 88990 31178 88998 31578
rect 88678 31168 88998 31178
rect 85684 29746 85694 30130
rect 86078 29746 86084 30130
rect 85684 25508 86084 29746
rect 89456 30130 89856 34368
rect 93228 34752 93628 38990
rect 97000 39374 97400 39600
rect 97000 38990 97010 39374
rect 97394 38990 97400 39374
rect 96284 36210 96484 38090
rect 96222 36200 96542 36210
rect 96222 35800 96234 36200
rect 96534 35800 96542 36200
rect 96222 35790 96542 35800
rect 93228 34368 93238 34752
rect 93622 34368 93628 34752
rect 92512 31588 92712 33468
rect 92450 31578 92770 31588
rect 92450 31178 92462 31578
rect 92762 31178 92770 31578
rect 92450 31168 92770 31178
rect 89456 29746 89466 30130
rect 89850 29746 89856 30130
rect 88740 26966 88940 28846
rect 88678 26956 88998 26966
rect 88678 26556 88690 26956
rect 88990 26556 88998 26956
rect 88678 26546 88998 26556
rect 85684 25124 85694 25508
rect 86078 25124 86084 25508
rect 85684 20886 86084 25124
rect 89456 25508 89856 29746
rect 93228 30130 93628 34368
rect 97000 34752 97400 38990
rect 97000 34368 97010 34752
rect 97394 34368 97400 34752
rect 96284 31588 96484 33468
rect 96222 31578 96542 31588
rect 96222 31178 96234 31578
rect 96534 31178 96542 31578
rect 96222 31168 96542 31178
rect 93228 29746 93238 30130
rect 93622 29746 93628 30130
rect 92512 26966 92712 28846
rect 92450 26956 92770 26966
rect 92450 26556 92462 26956
rect 92762 26556 92770 26956
rect 92450 26546 92770 26556
rect 89456 25124 89466 25508
rect 89850 25124 89856 25508
rect 88740 22344 88940 24224
rect 88678 22334 88998 22344
rect 88678 21934 88690 22334
rect 88990 21934 88998 22334
rect 88678 21924 88998 21934
rect 85684 20502 85694 20886
rect 86078 20502 86084 20886
rect 85684 16264 86084 20502
rect 89456 20886 89856 25124
rect 93228 25508 93628 29746
rect 97000 30130 97400 34368
rect 97000 29746 97010 30130
rect 97394 29746 97400 30130
rect 96284 26966 96484 28846
rect 96222 26956 96542 26966
rect 96222 26556 96234 26956
rect 96534 26556 96542 26956
rect 96222 26546 96542 26556
rect 93228 25124 93238 25508
rect 93622 25124 93628 25508
rect 92512 22344 92712 24224
rect 92450 22334 92770 22344
rect 92450 21934 92462 22334
rect 92762 21934 92770 22334
rect 92450 21924 92770 21934
rect 89456 20502 89466 20886
rect 89850 20502 89856 20886
rect 88740 17722 88940 19602
rect 88678 17712 88998 17722
rect 88678 17312 88690 17712
rect 88990 17312 88998 17712
rect 88678 17302 88998 17312
rect 85684 15880 85694 16264
rect 86078 15880 86084 16264
rect 85684 15000 86084 15880
rect 89456 16264 89856 20502
rect 93228 20886 93628 25124
rect 97000 25508 97400 29746
rect 97000 25124 97010 25508
rect 97394 25124 97400 25508
rect 96284 22344 96484 24224
rect 96222 22334 96542 22344
rect 96222 21934 96234 22334
rect 96534 21934 96542 22334
rect 96222 21924 96542 21934
rect 93228 20502 93238 20886
rect 93622 20502 93628 20886
rect 92512 17722 92712 19602
rect 92450 17712 92770 17722
rect 92450 17312 92462 17712
rect 92762 17312 92770 17712
rect 92450 17302 92770 17312
rect 89456 15880 89466 16264
rect 89850 15880 89856 16264
rect 89456 15000 89856 15880
rect 93228 16264 93628 20502
rect 97000 20886 97400 25124
rect 97000 20502 97010 20886
rect 97394 20502 97400 20886
rect 96284 17722 96484 19602
rect 96222 17712 96542 17722
rect 96222 17312 96234 17712
rect 96534 17312 96542 17712
rect 96222 17302 96542 17312
rect 93228 15880 93238 16264
rect 93622 15880 93628 16264
rect 93228 15000 93628 15880
rect 97000 16264 97400 20502
rect 97000 15880 97010 16264
rect 97394 15880 97400 16264
rect 97000 15000 97400 15880
rect 62336 13100 62536 14980
rect 66108 13100 66308 14980
rect 62274 13090 62594 13100
rect 62274 12690 62286 13090
rect 62586 12690 62594 13090
rect 62274 12680 62594 12690
rect 66046 13090 66366 13100
rect 66046 12690 66058 13090
rect 66358 12690 66366 13090
rect 66046 12680 66366 12690
rect 69880 12506 70080 14980
rect 88740 13100 88940 14980
rect 92512 13100 92712 14980
rect 96284 13100 96484 14980
rect 88678 13090 88998 13100
rect 88678 12690 88690 13090
rect 88990 12690 88998 13090
rect 88678 12680 88998 12690
rect 92450 13090 92770 13100
rect 92450 12690 92462 13090
rect 92762 12690 92770 13090
rect 92450 12680 92770 12690
rect 96222 13090 96542 13100
rect 96222 12690 96234 13090
rect 96534 12690 96542 13090
rect 96222 12680 96542 12690
rect 69818 12496 70138 12506
rect 69818 12096 69830 12496
rect 70130 12096 70138 12496
rect 69818 12086 70138 12096
rect 51730 5190 52136 5200
rect 52330 6610 52736 6620
rect 52330 6230 52340 6610
rect 52720 6410 52736 6610
rect 52720 6230 52730 6410
rect 51730 4810 51740 5190
rect 52120 4810 52130 5190
rect 51730 4800 52130 4810
rect 52330 4800 52730 6230
rect 40420 4550 40820 4560
rect 38620 4410 38870 4420
rect 37410 3870 37420 4250
rect 37790 3870 37800 4250
rect 37410 3860 37800 3870
rect 36640 3340 36650 3720
rect 37040 3340 37050 3720
rect 36640 2470 37050 3340
rect 38310 2700 38540 3300
rect 38220 2690 38620 2700
rect 38220 2310 38230 2690
rect 38610 2310 38620 2690
rect 38220 2300 38620 2310
rect 32870 1610 32880 1990
rect 33270 1610 33280 1990
rect 32870 1600 33280 1610
rect 38310 1480 38540 2300
rect 38220 1470 38620 1480
rect 38220 1090 38230 1470
rect 38610 1090 38620 1470
rect 38220 1080 38620 1090
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 200
rect 23370 0 23550 200
rect 27234 0 27414 200
use mosbius_col6 *mosbius_col6_0
timestamp 1757215509
transform 1 0 64370 0 1 35332
box -146 -32354 3794 8020
use mosbius_col6 *mosbius_col6_1
timestamp 1757215509
transform 1 0 68142 0 1 35332
box -146 -32354 3794 8020
use mosbius_col7 *mosbius_col7_0
timestamp 1757215509
transform 1 0 7790 0 1 35332
box -146 -32354 3794 8020
use mosbius_col7 *mosbius_col7_1
timestamp 1757215509
transform 1 0 11562 0 1 35332
box -146 -32354 3794 8020
use mosbius_col7 *mosbius_col7_2
timestamp 1757215509
transform 1 0 87002 0 1 35332
box -146 -32354 3794 8020
use mosbius_col7 *mosbius_col7_3
timestamp 1757215509
transform 1 0 83230 0 1 35332
box -146 -32354 3794 8020
use mosbius_col7 *mosbius_col7_4
timestamp 1757215509
transform 1 0 37966 0 1 35332
box -146 -32354 3794 8020
use mosbius_col7 *mosbius_col7_5
timestamp 1757215509
transform 1 0 41738 0 1 35332
box -146 -32354 3794 8020
use mosbius_col7 *mosbius_col7_6
timestamp 1757215509
transform 1 0 49282 0 1 35332
box -146 -32354 3794 8020
use mosbius_col7 *mosbius_col7_7
timestamp 1757215509
transform 1 0 45510 0 1 35332
box -146 -32354 3794 8020
use mosbius_col7 *mosbius_col7_8
timestamp 1757215509
transform 1 0 71914 0 1 35332
box -146 -32354 3794 8020
use mosbius_col8 *mosbius_col8_0
timestamp 1757215509
transform 1 0 4018 0 1 35332
box -146 -32354 3794 8020
use mosbius_col8 *mosbius_col8_1
timestamp 1757215509
transform 1 0 246 0 1 35332
box -146 -32354 3794 8020
use mosbius_col8 *mosbius_col8_2
timestamp 1757215509
transform 1 0 34194 0 1 35332
box -146 -32354 3794 8020
use mosbius_col8 *mosbius_col8_5
timestamp 1757215509
transform 1 0 15334 0 1 35332
box -146 -32354 3794 8020
use mosbius_col8 *mosbius_col8_6
timestamp 1757215509
transform 1 0 19106 0 1 35332
box -146 -32354 3794 8020
use mosbius_col8 *mosbius_col8_7
timestamp 1757215509
transform 1 0 22878 0 1 35332
box -146 -32354 3794 8020
use mosbius_col8 *mosbius_col8_8
timestamp 1757215509
transform 1 0 26650 0 1 35332
box -146 -32354 3794 8020
use mosbius_col8 *mosbius_col8_9
timestamp 1757215509
transform 1 0 30422 0 1 35332
box -146 -32354 3794 8020
use mosbius_col8 *mosbius_col8_10
timestamp 1757215509
transform 1 0 75686 0 1 35332
box -146 -32354 3794 8020
use mosbius_col8 *mosbius_col8_15
timestamp 1757215509
transform 1 0 53054 0 1 35332
box -146 -32354 3794 8020
use mosbius_col8 *mosbius_col8_16
timestamp 1757215509
transform 1 0 56826 0 1 35332
box -146 -32354 3794 8020
use mosbius_col8 *mosbius_col8_17
timestamp 1757215509
transform 1 0 60598 0 1 35332
box -146 -32354 3794 8020
use mosbius_col8 *mosbius_col8_22
timestamp 1757215509
transform 1 0 79458 0 1 35332
box -146 -32354 3794 8020
use mosbius_col8 *mosbius_col8_23
timestamp 1757215509
transform 1 0 90774 0 1 35332
box -146 -32354 3794 8020
use mosbius_col8 *mosbius_col8_25
timestamp 1757215509
transform 1 0 94546 0 1 35332
box -146 -32354 3794 8020
use sky130_fd_pr__nfet_g5v0d10v5_8ML6AG  sky130_fd_pr__nfet_g5v0d10v5_8ML6AG_0
timestamp 1757201930
transform 1 0 40671 0 1 5608
box -1621 -758 1621 758
use sky130_fd_pr__nfet_g5v0d10v5_8ML6AG  sky130_fd_pr__nfet_g5v0d10v5_8ML6AG_1
timestamp 1757201930
transform 1 0 49071 0 1 5608
box -1621 -758 1621 758
use sky130_fd_pr__nfet_g5v0d10v5_8263FJ *sky130_fd_pr__nfet_g5v0d10v5_8263FJ_1
timestamp 1757201930
transform -1 0 9573 0 -1 4967
box -673 -1367 673 1367
use sky130_fd_pr__nfet_g5v0d10v5_8263FJ *sky130_fd_pr__nfet_g5v0d10v5_8263FJ_2
timestamp 1757201930
transform -1 0 13273 0 -1 4967
box -673 -1367 673 1367
use sky130_fd_pr__nfet_g5v0d10v5_CLGMFJ  sky130_fd_pr__nfet_g5v0d10v5_CLGMFJ_0
timestamp 1757215441
transform 1 0 42411 0 1 2167
box -3811 -1367 3811 1367
use sky130_fd_pr__pfet_g5v0d10v5_AA5R3U  sky130_fd_pr__pfet_g5v0d10v5_AA5R3U_0
timestamp 1757201930
transform 1 0 68183 0 1 10315
box -2283 -1415 2283 1415
use sky130_fd_pr__pfet_g5v0d10v5_FGL9HY  sky130_fd_pr__pfet_g5v0d10v5_FGL9HY_0
timestamp 1757215542
transform 1 0 88985 0 1 2405
box -1335 -1415 1335 1415
use sky130_fd_pr__pfet_g5v0d10v5_FGL9HY  sky130_fd_pr__pfet_g5v0d10v5_FGL9HY_1
timestamp 1757215542
transform 1 0 88995 0 1 5725
box -1335 -1415 1335 1415
use sky130_fd_pr__pfet_g5v0d10v5_N4SDRF  sky130_fd_pr__pfet_g5v0d10v5_N4SDRF_0
timestamp 1757201930
transform -1 0 70241 0 -1 4551
box -3841 -2651 3841 2651
use sky130_fd_pr__pfet_g5v0d10v5_R4AJ4P  sky130_fd_pr__pfet_g5v0d10v5_R4AJ4P_0
timestamp 1757201930
transform 1 0 48735 0 1 2115
box -2035 -1415 2035 1415
<< labels >>
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 98624 45152
<< end >>
