magic
tech sky130A
magscale 1 2
timestamp 1757702553
<< viali >>
rect 1246 4228 3444 4262
rect 3410 2876 3444 4228
rect 1246 2842 3444 2876
rect 268 2532 3414 2566
rect 3380 162 3414 2532
rect 268 128 3414 162
<< metal1 >>
rect 888 4334 894 4340
rect 322 4300 894 4334
rect 82 4224 266 4230
rect 322 4208 356 4300
rect 402 4224 470 4230
rect 82 4164 266 4170
rect 402 4164 470 4170
rect 48 2842 82 4090
rect 520 3938 554 4300
rect 888 4288 894 4300
rect 946 4288 952 4340
rect 1060 4262 3456 4268
rect 1060 4228 1246 4262
rect 598 4170 604 4224
rect 672 4220 678 4224
rect 1060 4222 3410 4228
rect 1060 4220 1106 4222
rect 672 4174 1106 4220
rect 672 4170 678 4174
rect 272 3904 554 3938
rect 1282 4084 3260 4130
rect 272 3848 306 3904
rect 1282 3635 1328 4084
rect 652 3585 1328 3635
rect 652 3009 872 3059
rect 48 2796 176 2842
rect 826 2734 872 3009
rect 1282 3020 1328 3585
rect 1370 4046 1424 4052
rect 1370 3052 1424 3658
rect 1528 3446 1582 4052
rect 1528 3052 1582 3058
rect 1686 4046 1740 4052
rect 1686 3052 1740 3658
rect 1844 3446 1898 4052
rect 1844 3052 1898 3058
rect 2002 4046 2056 4052
rect 2002 3052 2056 3658
rect 2160 3446 2214 4052
rect 2160 3052 2214 3058
rect 2318 4046 2372 4052
rect 2318 3052 2372 3658
rect 2476 3446 2530 4052
rect 2476 3052 2530 3058
rect 2634 4046 2688 4052
rect 2634 3052 2688 3658
rect 2792 3446 2846 4052
rect 2792 3052 2846 3058
rect 2950 4046 3004 4052
rect 2950 3052 3004 3658
rect 3108 3446 3162 4052
rect 3108 3052 3162 3058
rect 3266 4046 3320 4052
rect 3266 3052 3320 3658
rect 1282 2974 3260 3020
rect 3398 2882 3410 4222
rect 1234 2876 3410 2882
rect 1234 2842 1246 2876
rect 3444 2842 3456 4262
rect 1234 2836 3456 2842
rect 164 2688 872 2734
rect 164 2434 210 2688
rect 662 2576 898 2582
rect 256 2566 662 2572
rect 898 2566 3426 2572
rect 256 2532 268 2566
rect 256 2526 662 2532
rect 898 2526 3380 2532
rect 662 2516 898 2522
rect 164 2388 3230 2434
rect 304 306 350 2388
rect 392 1808 446 2348
rect 392 740 446 1420
rect 392 346 446 352
rect 550 2342 604 2348
rect 550 1274 604 1954
rect 550 346 604 886
rect 708 1808 762 2348
rect 708 740 762 1420
rect 708 346 762 352
rect 866 2342 920 2348
rect 866 1274 920 1954
rect 866 346 920 886
rect 1024 1808 1078 2348
rect 1024 740 1078 1420
rect 1024 346 1078 352
rect 1182 2342 1236 2348
rect 1182 1274 1236 1954
rect 1182 346 1236 886
rect 1340 1808 1394 2348
rect 1340 740 1394 1420
rect 1340 346 1394 352
rect 1498 2342 1552 2348
rect 1498 1274 1552 1954
rect 1498 346 1552 886
rect 1656 1808 1710 2348
rect 1656 740 1710 1420
rect 1656 346 1710 352
rect 1814 2342 1868 2348
rect 1814 1274 1868 1954
rect 1814 346 1868 886
rect 1972 1808 2026 2348
rect 1972 740 2026 1420
rect 1972 346 2026 352
rect 2130 2342 2184 2348
rect 2130 1274 2184 1954
rect 2130 346 2184 886
rect 2288 1808 2342 2348
rect 2288 740 2342 1420
rect 2288 346 2342 352
rect 2446 2342 2500 2348
rect 2446 1274 2500 1954
rect 2446 346 2500 886
rect 2604 1808 2658 2348
rect 2604 740 2658 1420
rect 2604 346 2658 352
rect 2762 2342 2816 2348
rect 2762 1274 2816 1954
rect 2762 346 2816 886
rect 2920 1808 2974 2348
rect 2920 740 2974 1420
rect 2920 346 2974 352
rect 3078 2342 3132 2348
rect 3078 1274 3132 1954
rect 3078 346 3132 886
rect 3236 1808 3290 2348
rect 3236 740 3290 1420
rect 3236 346 3290 352
rect 304 260 3230 306
rect 3368 168 3380 2526
rect 256 162 3380 168
rect 256 128 268 162
rect 3414 128 3426 2566
rect 256 122 3426 128
<< via1 >>
rect 82 4170 266 4224
rect 402 4170 470 4224
rect 894 4288 946 4340
rect 604 4170 672 4224
rect 406 3694 498 3854
rect 448 3240 810 3404
rect 406 2790 498 2950
rect 1370 3658 1424 4046
rect 1528 3058 1582 3446
rect 1686 3658 1740 4046
rect 1844 3058 1898 3446
rect 2002 3658 2056 4046
rect 2160 3058 2214 3446
rect 2318 3658 2372 4046
rect 2476 3058 2530 3446
rect 2634 3658 2688 4046
rect 2792 3058 2846 3446
rect 2950 3658 3004 4046
rect 3108 3058 3162 3446
rect 3266 3658 3320 4046
rect 662 2566 898 2576
rect 662 2532 898 2566
rect 662 2522 898 2532
rect 392 1420 446 1808
rect 392 352 446 740
rect 550 1954 604 2342
rect 550 886 604 1274
rect 708 1420 762 1808
rect 708 352 762 740
rect 866 1954 920 2342
rect 866 886 920 1274
rect 1024 1420 1078 1808
rect 1024 352 1078 740
rect 1182 1954 1236 2342
rect 1182 886 1236 1274
rect 1340 1420 1394 1808
rect 1340 352 1394 740
rect 1498 1954 1552 2342
rect 1498 886 1552 1274
rect 1656 1420 1710 1808
rect 1656 352 1710 740
rect 1814 1954 1868 2342
rect 1814 886 1868 1274
rect 1972 1420 2026 1808
rect 1972 352 2026 740
rect 2130 1954 2184 2342
rect 2130 886 2184 1274
rect 2288 1420 2342 1808
rect 2288 352 2342 740
rect 2446 1954 2500 2342
rect 2446 886 2500 1274
rect 2604 1420 2658 1808
rect 2604 352 2658 740
rect 2762 1954 2816 2342
rect 2762 886 2816 1274
rect 2920 1420 2974 1808
rect 2920 352 2974 740
rect 3078 1954 3132 2342
rect 3078 886 3132 1274
rect 3236 1420 3290 1808
rect 3236 352 3290 740
<< metal2 >>
rect 882 4286 892 4342
rect 948 4286 958 4342
rect 82 4226 266 4230
rect 82 4224 92 4226
rect 256 4224 266 4226
rect 82 4168 92 4170
rect 256 4168 266 4170
rect 82 4164 266 4168
rect 398 4226 474 4230
rect 398 4224 408 4226
rect 464 4224 474 4226
rect 398 4170 402 4224
rect 470 4170 474 4224
rect 398 4168 408 4170
rect 464 4168 474 4170
rect 398 4164 474 4168
rect 600 4226 676 4230
rect 600 4224 610 4226
rect 666 4224 676 4226
rect 600 4170 604 4224
rect 672 4170 676 4224
rect 600 4168 610 4170
rect 666 4168 676 4170
rect 600 4164 676 4168
rect 1370 4046 3320 4052
rect 400 3694 406 3854
rect 498 3694 504 3854
rect 1370 3652 3320 3658
rect 1528 3446 3162 3452
rect 448 3404 810 3410
rect 448 3234 810 3240
rect 3002 3058 3108 3446
rect 1528 3052 3162 3058
rect 400 2790 406 2950
rect 498 2790 504 2950
rect 662 2580 898 2582
rect 662 2576 672 2580
rect 888 2576 898 2580
rect 662 2518 672 2522
rect 888 2518 898 2522
rect 662 2516 898 2518
rect 0 2342 3132 2348
rect 0 1954 10 2342
rect 0 1948 3132 1954
rect 3212 2338 3612 2348
rect 0 1280 292 1948
rect 3212 1824 3218 2338
rect 3606 1824 3612 2338
rect 3212 1814 3612 1824
rect 392 1808 3612 1814
rect 446 1420 708 1808
rect 762 1420 1024 1808
rect 1078 1420 1340 1808
rect 1394 1420 1656 1808
rect 1710 1420 1972 1808
rect 2026 1420 2288 1808
rect 2342 1420 2604 1808
rect 2658 1420 2920 1808
rect 2974 1420 3236 1808
rect 3290 1420 3612 1808
rect 392 1414 3612 1420
rect 0 1274 3132 1280
rect 0 886 550 1274
rect 604 886 866 1274
rect 920 886 1182 1274
rect 1236 886 1498 1274
rect 1552 886 1814 1274
rect 1868 886 2130 1274
rect 2184 886 2446 1274
rect 2500 886 2762 1274
rect 2816 886 3078 1274
rect 0 880 3132 886
rect 3212 746 3612 1414
rect 392 740 3612 746
rect 446 352 708 740
rect 762 352 1024 740
rect 1078 352 1340 740
rect 1394 352 1656 740
rect 1710 352 1972 740
rect 2026 352 2288 740
rect 2342 352 2604 740
rect 2658 352 2920 740
rect 2974 352 3236 740
rect 3290 352 3612 740
rect 392 346 3612 352
<< via2 >>
rect 892 4340 948 4342
rect 892 4288 894 4340
rect 894 4288 946 4340
rect 946 4288 948 4340
rect 892 4286 948 4288
rect 92 4224 256 4226
rect 92 4170 256 4224
rect 92 4168 256 4170
rect 408 4224 464 4226
rect 408 4170 464 4224
rect 408 4168 464 4170
rect 610 4224 666 4226
rect 610 4170 666 4224
rect 610 4168 666 4170
rect 406 3704 498 3844
rect 1380 3658 1424 4046
rect 1424 3658 1686 4046
rect 1686 3658 1740 4046
rect 1740 3658 2002 4046
rect 2002 3658 2056 4046
rect 2056 3658 2318 4046
rect 2318 3658 2372 4046
rect 2372 3658 2634 4046
rect 2634 3658 2688 4046
rect 2688 3658 2950 4046
rect 2950 3658 3004 4046
rect 3004 3658 3266 4046
rect 3266 3658 3310 4046
rect 458 3240 800 3404
rect 1538 3058 1582 3446
rect 1582 3058 1844 3446
rect 1844 3058 1898 3446
rect 1898 3058 2160 3446
rect 2160 3058 2214 3446
rect 2214 3058 2476 3446
rect 2476 3058 2530 3446
rect 2530 3058 2792 3446
rect 2792 3058 2846 3446
rect 2846 3058 3002 3446
rect 406 2800 498 2940
rect 672 2576 888 2580
rect 672 2522 888 2576
rect 672 2518 888 2522
rect 10 1954 550 2342
rect 550 1954 604 2342
rect 604 1954 866 2342
rect 866 1954 920 2342
rect 920 1954 1182 2342
rect 1182 1954 1236 2342
rect 1236 1954 1498 2342
rect 1498 1954 1552 2342
rect 1552 1954 1814 2342
rect 1814 1954 1868 2342
rect 1868 1954 2130 2342
rect 2130 1954 2184 2342
rect 2184 1954 2446 2342
rect 2446 1954 2500 2342
rect 2500 1954 2762 2342
rect 2762 1954 2816 2342
rect 2816 1954 3078 2342
rect 3078 1954 3122 2342
rect 3218 1824 3606 2338
<< metal3 >>
rect 886 4342 954 4352
rect 886 4286 892 4342
rect 948 4286 954 4342
rect 886 4276 954 4286
rect 20 4162 26 4232
rect 254 4226 262 4232
rect 256 4168 262 4226
rect 254 4162 262 4168
rect 340 4162 346 4232
rect 574 4226 672 4232
rect 574 4168 610 4226
rect 666 4168 672 4226
rect 890 4172 950 4276
rect 574 4162 672 4168
rect 1370 4050 3612 4052
rect 1370 4046 1752 4050
rect 1928 4046 3612 4050
rect 340 3694 346 3854
rect 574 3694 580 3854
rect 1370 3658 1380 4046
rect 3310 3658 3612 4046
rect 1370 3654 1752 3658
rect 1928 3654 3612 3658
rect 1370 3652 3612 3654
rect 1528 3446 3012 3452
rect 448 3404 666 3410
rect 448 3240 458 3404
rect 448 3234 666 3240
rect 894 3234 900 3410
rect 1528 3058 1538 3446
rect 3002 3058 3012 3446
rect 1528 3052 3012 3058
rect 340 2790 346 2950
rect 574 2790 580 2950
rect 1640 2750 2040 3052
rect 662 2582 898 2588
rect 662 2510 898 2516
rect 1640 2354 1752 2750
rect 1928 2354 2040 2750
rect 1640 2348 2040 2354
rect 0 2342 3132 2348
rect 0 1954 10 2342
rect 3122 1954 3132 2342
rect 0 1948 3132 1954
rect 3212 2338 3612 3652
rect 3212 1824 3218 2338
rect 3606 1824 3612 2338
rect 3212 1814 3612 1824
<< via3 >>
rect 26 4226 254 4232
rect 26 4168 92 4226
rect 92 4168 254 4226
rect 26 4162 254 4168
rect 346 4226 574 4232
rect 346 4168 408 4226
rect 408 4168 464 4226
rect 464 4168 574 4226
rect 346 4162 574 4168
rect 1752 4046 1928 4050
rect 346 3844 574 3854
rect 346 3704 406 3844
rect 406 3704 498 3844
rect 498 3704 574 3844
rect 346 3694 574 3704
rect 1752 3658 1928 4046
rect 1752 3654 1928 3658
rect 666 3404 894 3410
rect 666 3240 800 3404
rect 800 3240 894 3404
rect 666 3234 894 3240
rect 346 2940 574 2950
rect 346 2800 406 2940
rect 406 2800 498 2940
rect 498 2800 574 2940
rect 346 2790 574 2800
rect 662 2580 898 2582
rect 662 2518 672 2580
rect 672 2518 888 2580
rect 888 2518 898 2580
rect 662 2516 898 2518
rect 1752 2354 1928 2750
<< metal4 >>
rect 20 4232 260 4352
rect 20 4162 26 4232
rect 254 4162 260 4232
rect 20 0 260 4162
rect 340 4232 580 4352
rect 340 4162 346 4232
rect 574 4162 580 4232
rect 340 3854 580 4162
rect 340 3694 346 3854
rect 574 3694 580 3854
rect 340 2950 580 3694
rect 340 2790 346 2950
rect 574 2790 580 2950
rect 340 0 580 2790
rect 660 3410 900 4352
rect 1750 4050 1930 4352
rect 1750 3654 1752 4050
rect 1928 3654 1930 4050
rect 1750 3652 1930 3654
rect 660 3234 666 3410
rect 894 3234 900 3410
rect 660 2582 900 3234
rect 660 2516 662 2582
rect 898 2516 900 2582
rect 660 0 900 2516
rect 1750 2750 1930 2752
rect 1750 2354 1752 2750
rect 1928 2354 1930 2750
rect 1750 2352 1930 2354
use sky130_fd_pr__nfet_g5v0d10v5_SFRJCA  sky130_fd_pr__nfet_g5v0d10v5_SFRJCA_0
timestamp 1757702553
transform 1 0 2345 0 1 3552
box -1147 -758 1147 758
use sky130_fd_pr__pfet_g5v0d10v5_CYUY46  sky130_fd_pr__pfet_g5v0d10v5_CYUY46_0
timestamp 1757702553
transform 1 0 1841 0 1 1347
box -1651 -1297 1651 1297
use tt_lvl_shift  tt_lvl_shift_0
timestamp 1757702553
transform -1 0 880 0 -1 3322
box -2 -550 804 550
use tt_small_inv  tt_small_inv_0
timestamp 1757702553
transform 0 1 -4806 -1 0 4940
box 668 4844 940 5328
<< labels >>
rlabel metal4 20 0 260 4352 1 VDPWR
port 2 n power input
rlabel metal3 890 4172 950 4352 1 ctrl
port 4 n signal input
rlabel metal4 1750 3952 1930 4352 1 mod
port 5 n analog bidirectional
rlabel metal4 1750 2352 1930 2752 1 bus
port 6 n analog bidirectional
rlabel metal4 660 0 900 4352 1 VAPWR
port 3 n power input
rlabel metal4 340 0 580 4352 1 VGND
port 1 n ground input
<< properties >>
string FIXED_BBOX 0 0 3680 4352
<< end >>
