magic
tech sky130A
magscale 1 2
timestamp 1757298312
<< dnwell >>
rect 8500 4200 10700 7700
rect 12200 4200 14400 7700
rect 38700 5500 42700 7750
rect 47100 5500 51100 7750
<< nwell >>
rect 8420 7494 10780 7780
rect 8420 4406 8706 7494
rect 10494 4406 10780 7494
rect 8420 4120 10780 4406
rect 12120 7494 14480 7780
rect 12120 4406 12406 7494
rect 14194 4406 14480 7494
rect 38620 7544 42780 7830
rect 38620 5706 38906 7544
rect 42494 5706 42780 7544
rect 38620 5420 42780 5706
rect 47020 7544 51180 7830
rect 47020 5706 47306 7544
rect 50894 5706 51180 7544
rect 47020 5420 51180 5706
rect 12120 4120 14480 4406
<< nsubdiff >>
rect 38657 7773 42743 7793
rect 8457 7723 10743 7743
rect 8457 7689 8537 7723
rect 10663 7689 10743 7723
rect 8457 7669 10743 7689
rect 8457 7663 8531 7669
rect 8457 4237 8477 7663
rect 8511 4237 8531 7663
rect 8457 4231 8531 4237
rect 10669 7663 10743 7669
rect 10669 4237 10689 7663
rect 10723 4237 10743 7663
rect 10669 4231 10743 4237
rect 8457 4211 10743 4231
rect 8457 4177 8537 4211
rect 10663 4177 10743 4211
rect 8457 4157 10743 4177
rect 12157 7723 14443 7743
rect 12157 7689 12237 7723
rect 14363 7689 14443 7723
rect 12157 7669 14443 7689
rect 12157 7663 12231 7669
rect 12157 4237 12177 7663
rect 12211 4237 12231 7663
rect 12157 4231 12231 4237
rect 14369 7663 14443 7669
rect 14369 4237 14389 7663
rect 14423 4237 14443 7663
rect 38657 7739 38737 7773
rect 42663 7739 42743 7773
rect 38657 7719 42743 7739
rect 38657 7713 38731 7719
rect 38657 5537 38677 7713
rect 38711 5537 38731 7713
rect 38657 5531 38731 5537
rect 42669 7713 42743 7719
rect 42669 5537 42689 7713
rect 42723 5537 42743 7713
rect 42669 5531 42743 5537
rect 38657 5511 42743 5531
rect 38657 5477 38737 5511
rect 42663 5477 42743 5511
rect 38657 5457 42743 5477
rect 47057 7773 51143 7793
rect 47057 7739 47137 7773
rect 51063 7739 51143 7773
rect 47057 7719 51143 7739
rect 47057 7713 47131 7719
rect 47057 5537 47077 7713
rect 47111 5537 47131 7713
rect 47057 5531 47131 5537
rect 51069 7713 51143 7719
rect 51069 5537 51089 7713
rect 51123 5537 51143 7713
rect 51069 5531 51143 5537
rect 47057 5511 51143 5531
rect 47057 5477 47137 5511
rect 51063 5477 51143 5511
rect 47057 5457 51143 5477
rect 14369 4231 14443 4237
rect 12157 4211 14443 4231
rect 12157 4177 12237 4211
rect 14363 4177 14443 4211
rect 12157 4157 14443 4177
<< nsubdiffcont >>
rect 8537 7689 10663 7723
rect 8477 4237 8511 7663
rect 10689 4237 10723 7663
rect 8537 4177 10663 4211
rect 12237 7689 14363 7723
rect 12177 4237 12211 7663
rect 14389 4237 14423 7663
rect 38737 7739 42663 7773
rect 38677 5537 38711 7713
rect 42689 5537 42723 7713
rect 38737 5477 42663 5511
rect 47137 7739 51063 7773
rect 47077 5537 47111 7713
rect 51089 5537 51123 7713
rect 47137 5477 51063 5511
rect 12237 4177 14363 4211
<< locali >>
rect 26940 44620 27170 44630
rect 26756 44550 26874 44552
rect 26510 44540 26874 44550
rect 26510 44460 26520 44540
rect 26870 44460 26874 44540
rect 26510 44450 26874 44460
rect 26940 44450 26960 44620
rect 27160 44450 27170 44620
rect 26940 44440 27170 44450
rect 65660 12640 70700 13000
rect 65660 10000 66280 12640
rect 70090 10000 70700 12640
rect 65660 9640 70700 10000
rect 7900 8190 14900 8200
rect 7900 7710 8220 8190
rect 8900 7723 12010 8190
rect 12690 7723 14900 8190
rect 10663 7710 12010 7723
rect 7900 7689 8537 7710
rect 10663 7689 12237 7710
rect 14363 7689 14900 7723
rect 7900 7663 8511 7689
rect 7900 4237 8477 7663
rect 10689 7663 12211 7689
rect 8760 7260 10380 7460
rect 8760 7020 8960 7260
rect 10180 7040 10380 7260
rect 8760 6140 9100 7020
rect 10040 6160 10380 7040
rect 8760 5800 8960 6140
rect 10180 5800 10380 6160
rect 8760 4920 9100 5800
rect 10040 4920 10380 5800
rect 8760 4680 8960 4920
rect 10180 4680 10380 4920
rect 8760 4480 10380 4680
rect 7900 4211 8511 4237
rect 10723 4237 12177 7663
rect 14389 7663 14900 7689
rect 12460 7260 14080 7460
rect 12460 7020 12660 7260
rect 13880 7020 14080 7260
rect 12460 6140 12800 7020
rect 13740 6140 14080 7020
rect 12460 5800 12660 6140
rect 13880 5820 14080 6140
rect 12460 4920 12800 5800
rect 13740 4940 14080 5820
rect 12460 4680 12660 4920
rect 13880 4680 14080 4940
rect 12460 4480 14080 4680
rect 10689 4211 12211 4237
rect 14423 4237 14900 7663
rect 38290 7773 43100 8160
rect 66160 8100 74110 8390
rect 38290 7739 38737 7773
rect 42663 7739 43100 7773
rect 38290 7713 38711 7739
rect 38290 6040 38677 7713
rect 42689 7713 43100 7739
rect 39030 7290 42320 7590
rect 39030 7100 39400 7290
rect 41950 7100 42320 7290
rect 39030 6120 39410 7100
rect 41930 6120 42320 7100
rect 38711 6040 38870 6050
rect 38290 5420 38630 6040
rect 38860 5511 38870 6040
rect 39030 5920 39400 6120
rect 41950 5920 42320 6120
rect 39030 5620 42320 5920
rect 42723 5537 43100 7713
rect 46800 7773 51400 8070
rect 46800 7739 47137 7773
rect 51063 7739 51400 7773
rect 46800 7713 47111 7739
rect 46800 6800 47077 7713
rect 46730 6790 47077 6800
rect 51089 7713 51400 7739
rect 46730 6410 46740 6790
rect 46730 6400 47077 6410
rect 42689 5511 43100 5537
rect 42663 5477 43100 5511
rect 38860 5420 43100 5477
rect 38290 5100 43100 5420
rect 46800 5537 47077 6400
rect 47430 7290 50720 7590
rect 47430 7100 47800 7290
rect 50350 7100 50720 7290
rect 47430 6120 47810 7100
rect 50330 6120 50720 7100
rect 47430 5920 47800 6120
rect 50350 5920 50720 6120
rect 47430 5620 50720 5920
rect 46800 5511 47111 5537
rect 51123 5537 51400 7713
rect 51089 5511 51400 5537
rect 46800 5477 47137 5511
rect 51063 5477 51400 5511
rect 46800 5190 51400 5477
rect 14389 4211 14900 4237
rect 7900 4177 8537 4211
rect 10663 4177 12237 4211
rect 14363 4177 14900 4211
rect 7900 3700 14900 4177
rect 38460 4470 46350 4670
rect 38460 4260 39000 4470
rect 45830 4260 46350 4470
rect 38460 3300 39070 4260
rect 45760 3300 46350 4260
rect 38460 3050 39000 3300
rect 38460 2090 39070 3050
rect 45830 3040 46350 3300
rect 38460 1870 39000 2090
rect 45760 2080 46350 3040
rect 45840 1870 46350 2080
rect 38460 1670 46350 1870
rect 46780 4430 50690 4560
rect 46780 4230 47170 4430
rect 46780 3250 47200 4230
rect 50300 4220 50690 4430
rect 46780 2990 47170 3250
rect 50270 3240 50690 4220
rect 50300 2990 50690 3240
rect 46780 2010 47200 2990
rect 50270 2010 50690 2990
rect 66160 3010 66880 8100
rect 73600 3010 74110 8100
rect 83760 8050 86680 8280
rect 83760 5400 84260 8050
rect 86180 5400 86680 8050
rect 83760 5180 86680 5400
rect 66160 2650 74110 3010
rect 83760 4720 86660 4960
rect 46780 1800 47170 2010
rect 50300 1800 50690 2010
rect 83760 2100 84250 4720
rect 86170 2100 86660 4720
rect 83760 1860 86660 2100
rect 46780 1670 50690 1800
rect 51760 1190 52280 1250
rect 51760 1030 51930 1190
rect 51760 830 52050 1030
rect 51760 670 51930 830
rect 52230 670 52280 1190
rect 51760 590 52280 670
rect 52340 1120 52880 1250
rect 52340 740 52390 1120
rect 52700 970 52880 1120
rect 52570 960 52880 970
rect 52570 900 52680 960
rect 52830 900 52880 960
rect 52570 890 52880 900
rect 52700 740 52880 890
rect 52340 590 52880 740
<< viali >>
rect 26520 44460 26870 44540
rect 26960 44450 27160 44620
rect 8220 7723 8900 8190
rect 12010 7723 12690 8190
rect 8220 7710 8537 7723
rect 8537 7710 8900 7723
rect 12010 7710 12237 7723
rect 12237 7710 12690 7723
rect 38630 5537 38677 6040
rect 38677 5537 38711 6040
rect 38711 5537 38860 6040
rect 38630 5511 38860 5537
rect 46740 6410 47077 6790
rect 47077 6410 47100 6790
rect 38630 5477 38737 5511
rect 38737 5477 38860 5511
rect 38630 5420 38860 5477
rect 52680 900 52830 960
<< metal1 >>
rect 2990 45140 3090 45150
rect 2990 44840 3000 45140
rect 3080 44970 3090 45140
rect 3540 45140 3640 45150
rect 3540 44970 3550 45140
rect 3080 44840 3550 44970
rect 3630 44970 3640 45140
rect 4100 45140 4200 45150
rect 4100 44970 4110 45140
rect 3630 44840 4110 44970
rect 4190 44970 4200 45140
rect 4650 45140 4750 45150
rect 4650 44970 4660 45140
rect 4190 44840 4660 44970
rect 4740 44970 4750 45140
rect 5200 45140 5300 45150
rect 5200 44970 5210 45140
rect 4740 44840 5210 44970
rect 5290 44970 5300 45140
rect 5760 45140 5860 45150
rect 5760 44970 5770 45140
rect 5290 44840 5770 44970
rect 5850 44970 5860 45140
rect 6310 45140 6410 45150
rect 6310 44970 6320 45140
rect 5850 44840 6320 44970
rect 6400 44970 6410 45140
rect 6860 45140 6960 45150
rect 6860 44970 6870 45140
rect 6400 44840 6870 44970
rect 6950 44970 6960 45140
rect 7400 45140 7500 45150
rect 7400 44970 7410 45140
rect 6950 44840 7410 44970
rect 7490 44970 7500 45140
rect 7960 45140 8060 45150
rect 7960 44970 7970 45140
rect 7490 44840 7970 44970
rect 8050 44970 8060 45140
rect 8500 45140 8600 45150
rect 8500 44970 8510 45140
rect 8050 44840 8510 44970
rect 8590 44970 8600 45140
rect 9060 45140 9160 45150
rect 9060 44970 9070 45140
rect 8590 44840 9070 44970
rect 9150 44970 9160 45140
rect 9610 45140 9710 45150
rect 9610 44970 9620 45140
rect 9150 44840 9620 44970
rect 9700 44970 9710 45140
rect 10170 45140 10270 45150
rect 10170 44970 10180 45140
rect 9700 44840 10180 44970
rect 10260 44970 10270 45140
rect 10720 45140 10820 45150
rect 10720 44970 10730 45140
rect 10260 44840 10730 44970
rect 10810 44970 10820 45140
rect 11280 45140 11380 45150
rect 11280 44970 11290 45140
rect 10810 44840 11290 44970
rect 11370 44970 11380 45140
rect 12380 45140 12480 45150
rect 12380 44970 12390 45140
rect 11370 44960 12390 44970
rect 11370 44840 11890 44960
rect 2990 44830 11890 44840
rect 11880 44770 11890 44830
rect 12140 44840 12390 44960
rect 12470 44970 12480 45140
rect 12930 45140 13030 45150
rect 12930 44970 12940 45140
rect 12470 44840 12940 44970
rect 13020 44970 13030 45140
rect 13470 45140 13570 45150
rect 13470 44970 13480 45140
rect 13020 44840 13480 44970
rect 13560 44970 13570 45140
rect 14030 45140 14130 45150
rect 14030 44970 14040 45140
rect 13560 44840 14040 44970
rect 14120 44970 14130 45140
rect 14580 45140 14680 45150
rect 14580 44970 14590 45140
rect 14120 44840 14590 44970
rect 14670 44970 14680 45140
rect 15130 45140 15230 45150
rect 15130 44970 15140 45140
rect 14670 44840 15140 44970
rect 15220 44970 15230 45140
rect 16240 45140 16340 45150
rect 16240 44970 16250 45140
rect 15220 44840 16250 44970
rect 16330 44970 16340 45140
rect 16790 45140 16890 45150
rect 16790 44970 16800 45140
rect 16330 44840 16800 44970
rect 16880 44970 16890 45140
rect 17340 45140 17440 45150
rect 17340 44970 17350 45140
rect 16880 44840 17350 44970
rect 17430 44970 17440 45140
rect 17900 45140 18000 45150
rect 17900 44970 17910 45140
rect 17430 44840 17910 44970
rect 17990 44970 18000 45140
rect 18450 45140 18550 45150
rect 18450 44970 18460 45140
rect 17990 44840 18460 44970
rect 18540 44970 18550 45140
rect 19000 45140 19100 45150
rect 19000 44970 19010 45140
rect 18540 44840 19010 44970
rect 19090 44970 19100 45140
rect 19550 45140 19650 45150
rect 19550 44970 19560 45140
rect 19090 44840 19560 44970
rect 19640 44970 19650 45140
rect 20110 45140 20210 45150
rect 20110 44970 20120 45140
rect 19640 44840 20120 44970
rect 20200 44970 20210 45140
rect 20660 45140 20760 45150
rect 20660 44970 20670 45140
rect 20200 44840 20670 44970
rect 20750 44970 20760 45140
rect 21210 45140 21310 45150
rect 21210 44970 21220 45140
rect 20750 44840 21220 44970
rect 21300 44970 21310 45140
rect 21760 45140 21860 45150
rect 21760 44970 21770 45140
rect 21300 44840 21770 44970
rect 21850 44970 21860 45140
rect 22300 45140 22400 45150
rect 22300 44970 22310 45140
rect 21850 44840 22310 44970
rect 22390 44970 22400 45140
rect 23970 45140 24070 45150
rect 23970 44970 23980 45140
rect 22390 44840 23980 44970
rect 24060 44840 24070 45140
rect 12140 44830 24070 44840
rect 24470 45140 24660 45150
rect 24470 44960 24480 45140
rect 24650 44960 24660 45140
rect 12140 44770 12150 44830
rect 11880 44760 12150 44770
rect 3500 44580 3650 44590
rect 24470 44580 24660 44960
rect 3500 44440 3510 44580
rect 3640 44440 24660 44580
rect 25570 45140 25760 45150
rect 25570 44960 25580 45140
rect 25750 44960 25760 45140
rect 25570 44580 25760 44960
rect 27000 45010 27220 45020
rect 27000 44930 27010 45010
rect 26730 44870 27010 44930
rect 27210 44870 27220 45010
rect 26730 44660 27220 44870
rect 26940 44620 28370 44630
rect 25570 44540 26890 44580
rect 25570 44460 26520 44540
rect 26870 44460 26890 44540
rect 25570 44440 26890 44460
rect 26940 44450 26960 44620
rect 27160 44450 28110 44620
rect 28360 44450 28370 44620
rect 26940 44440 28370 44450
rect 3500 44430 3650 44440
rect 66230 12960 70990 12970
rect 66230 12770 70610 12960
rect 70980 12770 70990 12960
rect 66230 12760 70990 12770
rect 66320 12690 66570 12700
rect 66320 12500 66330 12690
rect 66560 12500 66570 12690
rect 66320 12480 66570 12500
rect 66640 12490 66890 12760
rect 66950 12690 67200 12700
rect 66950 12500 66960 12690
rect 67190 12500 67200 12690
rect 66950 12490 67200 12500
rect 66250 12420 66310 12430
rect 66250 11440 66310 11450
rect 66250 11180 66310 11190
rect 66250 10200 66310 10210
rect 66350 10150 66380 12480
rect 66420 12420 66480 12430
rect 66420 11440 66480 11450
rect 66420 11180 66480 11190
rect 66420 10200 66480 10210
rect 66510 10150 66540 12480
rect 66570 12420 66630 12430
rect 66570 11440 66630 11450
rect 66570 11180 66630 11190
rect 66570 10200 66630 10210
rect 66670 10150 66700 12490
rect 66730 12420 66790 12430
rect 66730 11440 66790 11450
rect 66730 11180 66790 11190
rect 66730 10200 66790 10210
rect 66830 10150 66860 12490
rect 66890 12420 66950 12430
rect 66890 11440 66950 11450
rect 66890 11180 66950 11190
rect 66890 10200 66950 10210
rect 66980 10150 67010 12490
rect 67050 12420 67110 12430
rect 67050 11440 67110 11450
rect 67050 11180 67110 11190
rect 67050 10200 67110 10210
rect 67140 10150 67170 12490
rect 67270 12480 67520 12760
rect 67590 12690 67840 12700
rect 67590 12500 67600 12690
rect 67830 12500 67840 12690
rect 67590 12490 67840 12500
rect 67200 12420 67260 12430
rect 67200 11440 67260 11450
rect 67200 11180 67260 11190
rect 67200 10200 67260 10210
rect 52930 10090 53290 10100
rect 52930 9490 53010 10090
rect 53280 9490 53290 10090
rect 66320 9870 66570 10150
rect 66640 10130 66880 10150
rect 66640 9940 66650 10130
rect 66870 9940 66880 10130
rect 66640 9930 66880 9940
rect 66960 9870 67200 10150
rect 67300 10140 67330 12480
rect 67360 12420 67420 12430
rect 67360 11440 67420 11450
rect 67360 11180 67420 11190
rect 67360 10200 67420 10210
rect 67460 10140 67490 12480
rect 67520 12420 67580 12430
rect 67520 11440 67580 11450
rect 67520 11180 67580 11190
rect 67520 10200 67580 10210
rect 67620 10150 67650 12490
rect 67680 12420 67740 12430
rect 67680 11440 67740 11450
rect 67680 11180 67740 11190
rect 67680 10200 67740 10210
rect 67770 10150 67800 12490
rect 67930 12480 68180 12760
rect 68220 12690 68470 12700
rect 68220 12500 68230 12690
rect 68460 12500 68470 12690
rect 68220 12490 68470 12500
rect 67840 12420 67900 12430
rect 67840 11440 67900 11450
rect 67840 11180 67900 11190
rect 67840 10200 67900 10210
rect 67270 10130 67520 10140
rect 67270 9940 67280 10130
rect 67510 9940 67520 10130
rect 67270 9930 67520 9940
rect 67590 9870 67840 10150
rect 67930 10140 67960 12480
rect 67990 12420 68050 12430
rect 67990 11440 68050 11450
rect 67990 11180 68050 11190
rect 67990 10200 68050 10210
rect 68090 10140 68120 12480
rect 68150 12420 68210 12430
rect 68150 11440 68210 11450
rect 68150 11180 68210 11190
rect 68150 10200 68210 10210
rect 68250 10150 68280 12490
rect 68310 12420 68370 12430
rect 68310 11440 68370 11450
rect 68310 11180 68370 11190
rect 68310 10200 68370 10210
rect 68410 10150 68440 12490
rect 68530 12480 68780 12760
rect 68850 12690 69100 12700
rect 68850 12500 68860 12690
rect 69090 12500 69100 12690
rect 68850 12490 69100 12500
rect 68470 12420 68530 12430
rect 68470 11440 68530 11450
rect 68470 11180 68530 11190
rect 68470 10200 68530 10210
rect 67900 10130 68150 10140
rect 67900 9940 67910 10130
rect 68140 9940 68150 10130
rect 67900 9930 68150 9940
rect 68220 9870 68470 10150
rect 68560 10140 68590 12480
rect 68630 12420 68690 12430
rect 68630 11440 68690 11450
rect 68630 11180 68690 11190
rect 68630 10200 68690 10210
rect 68720 10140 68750 12480
rect 68780 12420 68840 12430
rect 68780 11440 68840 11450
rect 68780 11180 68840 11190
rect 68780 10200 68840 10210
rect 68880 10150 68910 12490
rect 68940 12420 69000 12430
rect 68940 11440 69000 11450
rect 68940 11180 69000 11190
rect 68940 10200 69000 10210
rect 69040 10150 69070 12490
rect 69170 12480 69420 12760
rect 69480 12690 69730 12700
rect 69480 12500 69490 12690
rect 69720 12500 69730 12690
rect 69480 12490 69730 12500
rect 69100 12420 69160 12430
rect 69100 11440 69160 11450
rect 69100 11180 69160 11190
rect 69100 10200 69160 10210
rect 68530 10130 68780 10140
rect 68530 9940 68540 10130
rect 68770 9940 68780 10130
rect 68530 9930 68780 9940
rect 68850 9870 69100 10150
rect 69190 10140 69220 12480
rect 69260 12420 69320 12430
rect 69260 11440 69320 11450
rect 69260 11180 69320 11190
rect 69260 10200 69320 10210
rect 69350 10140 69380 12480
rect 69420 12420 69480 12430
rect 69420 11440 69480 11450
rect 69420 11180 69480 11190
rect 69420 10200 69480 10210
rect 69510 10150 69540 12490
rect 69580 12420 69640 12430
rect 69580 11440 69640 11450
rect 69580 11180 69640 11190
rect 69580 10200 69640 10210
rect 69670 10150 69700 12490
rect 69800 12480 70050 12760
rect 69730 12420 69790 12430
rect 69730 11440 69790 11450
rect 69730 11180 69790 11190
rect 69730 10200 69790 10210
rect 69170 10130 69410 10140
rect 69170 9940 69180 10130
rect 69400 9940 69410 10130
rect 69170 9930 69410 9940
rect 69480 9870 69730 10150
rect 69830 10140 69860 12480
rect 69890 12420 69950 12430
rect 69890 11440 69950 11450
rect 69890 11180 69950 11190
rect 69890 10200 69950 10210
rect 69990 10140 70020 12480
rect 70060 12420 70120 12430
rect 70060 11440 70120 11450
rect 70060 11180 70120 11190
rect 70060 10200 70120 10210
rect 69800 10130 70040 10140
rect 69800 9940 69810 10130
rect 70030 9940 70040 10130
rect 69800 9930 70040 9940
rect 66230 9860 71590 9870
rect 66230 9670 71210 9860
rect 71580 9670 71590 9860
rect 66230 9660 71590 9670
rect 52930 9480 53290 9490
rect 52930 8650 53230 9480
rect 71190 8910 71870 8920
rect 71190 8710 71200 8910
rect 71860 8710 71870 8910
rect 71190 8700 71870 8710
rect 8200 8190 8920 8200
rect 8200 7710 8220 8190
rect 8900 7710 8920 8190
rect 8200 7700 8920 7710
rect 11990 8190 12710 8200
rect 11990 7710 12010 8190
rect 12690 7710 12710 8190
rect 11990 7700 12710 7710
rect 13070 7200 13150 8580
rect 13390 7200 13470 8580
rect 52520 8400 53230 8650
rect 41180 8120 42520 8130
rect 41180 7840 41190 8120
rect 41560 7840 42210 8120
rect 42510 7840 42520 8120
rect 41180 7830 42520 7840
rect 39440 7410 45190 7420
rect 39440 7220 44800 7410
rect 8720 7120 10080 7200
rect 12780 7120 14100 7200
rect 8720 6040 8860 7120
rect 9880 7070 10040 7080
rect 9100 7060 9260 7070
rect 9100 6100 9110 7060
rect 9250 6100 9260 7060
rect 9100 6090 9260 6100
rect 9370 7060 9450 7070
rect 9370 6100 9380 7060
rect 9440 6100 9450 7060
rect 9370 6090 9450 6100
rect 9530 7060 9610 7070
rect 9530 6100 9540 7060
rect 9600 6100 9610 7060
rect 9530 6090 9610 6100
rect 9690 7060 9770 7070
rect 9690 6100 9700 7060
rect 9760 6100 9770 7060
rect 9880 6110 9890 7070
rect 10030 6110 10040 7070
rect 9880 6100 10040 6110
rect 12800 7060 12960 7070
rect 12800 6100 12810 7060
rect 12950 6100 12960 7060
rect 9690 6090 9770 6100
rect 12800 6090 12960 6100
rect 13070 7060 13150 7120
rect 13070 6100 13080 7060
rect 13140 6100 13150 7060
rect 13070 6090 13150 6100
rect 13230 7060 13310 7070
rect 13230 6100 13240 7060
rect 13300 6100 13310 7060
rect 13230 6090 13310 6100
rect 13390 7060 13470 7120
rect 13390 6100 13400 7060
rect 13460 6100 13470 7060
rect 13590 7060 13750 7070
rect 13590 7020 13600 7060
rect 13580 6140 13600 7020
rect 13390 6090 13470 6100
rect 13590 6100 13600 6140
rect 13740 6100 13750 7060
rect 13590 6090 13750 6100
rect 13960 6040 14100 7120
rect 39230 7100 39400 7190
rect 39460 7160 39510 7220
rect 39620 7160 39670 7220
rect 40090 7160 40140 7220
rect 40250 7160 40300 7220
rect 40720 7160 40770 7220
rect 40880 7160 40930 7220
rect 41350 7160 41400 7220
rect 41520 7160 41570 7220
rect 39230 7090 39420 7100
rect 39230 6130 39240 7090
rect 39410 6130 39420 7090
rect 39230 6120 39420 6130
rect 8720 5900 10080 6040
rect 12780 5900 14100 6040
rect 8720 5320 8860 5900
rect 8560 5310 8860 5320
rect 8560 5130 8570 5310
rect 8850 5130 8860 5310
rect 8560 5120 8860 5130
rect 8720 4820 8860 5120
rect 9100 5840 9260 5850
rect 9100 4880 9110 5840
rect 9250 4880 9260 5840
rect 9100 4870 9260 4880
rect 9370 5840 9450 5850
rect 9370 4880 9380 5840
rect 9440 4880 9450 5840
rect 9370 4870 9450 4880
rect 9530 5840 9610 5850
rect 9530 4880 9540 5840
rect 9600 4880 9610 5840
rect 9530 4870 9610 4880
rect 9690 5840 9770 5850
rect 9690 4880 9700 5840
rect 9760 4880 9770 5840
rect 9690 4870 9770 4880
rect 9880 5840 10040 5850
rect 9880 4880 9890 5840
rect 10030 4880 10040 5840
rect 9880 4870 10040 4880
rect 12800 5840 12960 5850
rect 12800 4880 12810 5840
rect 12950 4880 12960 5840
rect 12800 4870 12960 4880
rect 13070 5840 13150 5850
rect 13070 4880 13080 5840
rect 13140 4880 13150 5840
rect 13070 4870 13150 4880
rect 13230 5840 13310 5850
rect 13230 4880 13240 5840
rect 13300 4880 13310 5840
rect 13230 4870 13310 4880
rect 13390 5840 13470 5850
rect 13390 4880 13400 5840
rect 13460 4880 13470 5840
rect 13590 5840 13750 5850
rect 13590 5820 13600 5840
rect 13580 4940 13600 5820
rect 13390 4870 13470 4880
rect 13590 4880 13600 4940
rect 13740 4880 13750 5840
rect 13590 4870 13750 4880
rect 13960 5320 14100 5900
rect 38620 6040 38870 6060
rect 38620 5420 38630 6040
rect 38860 5420 38870 6040
rect 39230 6030 39400 6120
rect 39470 6050 39500 7160
rect 39540 7090 39600 7100
rect 39540 6120 39600 6130
rect 39630 6050 39660 7160
rect 39690 7090 39750 7100
rect 39690 6120 39750 6130
rect 39780 6050 39810 7160
rect 39850 7090 39910 7100
rect 39850 6120 39910 6130
rect 39940 6050 39970 7160
rect 40010 7090 40070 7100
rect 40010 6120 40070 6130
rect 40100 6050 40130 7160
rect 40170 7090 40230 7100
rect 40170 6120 40230 6130
rect 40260 6050 40290 7160
rect 40330 7090 40390 7100
rect 40330 6120 40390 6130
rect 40420 6050 40450 7160
rect 40480 7090 40540 7100
rect 40480 6120 40540 6130
rect 40580 6050 40610 7160
rect 40640 7090 40700 7100
rect 40640 6120 40700 6130
rect 40730 6050 40760 7160
rect 40800 7090 40860 7100
rect 40800 6120 40860 6130
rect 40890 6050 40920 7160
rect 40960 7090 41020 7100
rect 40960 6120 41020 6130
rect 41050 6050 41080 7160
rect 41120 7090 41180 7100
rect 41120 6120 41180 6130
rect 41210 6050 41240 7160
rect 41270 7090 41330 7100
rect 41270 6120 41330 6130
rect 41360 6050 41390 7160
rect 41430 7090 41490 7100
rect 41430 6120 41490 6130
rect 41530 6050 41560 7160
rect 41590 7090 41650 7100
rect 41590 6120 41650 6130
rect 41680 6050 41710 7160
rect 41750 7090 41810 7100
rect 41750 6120 41810 6130
rect 41850 6050 41880 7160
rect 41950 7100 42120 7190
rect 41930 7090 42120 7100
rect 41930 6130 41940 7090
rect 42110 6130 42120 7090
rect 44790 7030 44800 7220
rect 45180 7030 45190 7410
rect 47840 7410 51290 7420
rect 47840 7230 50730 7410
rect 51280 7230 51290 7410
rect 47840 7220 51290 7230
rect 44790 7020 45190 7030
rect 47560 7100 47800 7190
rect 47860 7160 47910 7220
rect 48020 7160 48070 7220
rect 48490 7160 48540 7220
rect 48650 7160 48700 7220
rect 49120 7160 49170 7220
rect 49280 7160 49330 7220
rect 49750 7160 49800 7220
rect 49920 7160 49970 7220
rect 47560 7090 47820 7100
rect 46720 6790 47120 6800
rect 46720 6410 46740 6790
rect 47100 6410 47120 6790
rect 46720 6400 47120 6410
rect 41930 6120 42120 6130
rect 39780 6000 39830 6050
rect 39930 6000 39980 6050
rect 40410 6000 40460 6050
rect 40570 6000 40620 6050
rect 41040 6000 41090 6050
rect 41200 6000 41250 6050
rect 41670 6000 41720 6050
rect 41840 6000 41890 6050
rect 41950 6030 42120 6120
rect 44190 6190 44590 6200
rect 44190 6000 44200 6190
rect 39440 5810 44200 6000
rect 44580 6000 44590 6190
rect 47560 6130 47640 7090
rect 47810 6130 47820 7090
rect 47560 6120 47820 6130
rect 44580 5810 45180 6000
rect 39440 5800 45180 5810
rect 38620 5400 38870 5420
rect 13960 5310 14260 5320
rect 13960 5130 13970 5310
rect 14250 5130 14260 5310
rect 47560 5290 47800 6120
rect 47870 6050 47900 7160
rect 47940 7090 48000 7100
rect 47940 6120 48000 6130
rect 48030 6050 48060 7160
rect 48090 7090 48150 7100
rect 48090 6120 48150 6130
rect 48180 6050 48210 7160
rect 48250 7090 48310 7100
rect 48250 6120 48310 6130
rect 48340 6050 48370 7160
rect 48410 7090 48470 7100
rect 48410 6120 48470 6130
rect 48500 6050 48530 7160
rect 48570 7090 48630 7100
rect 48570 6120 48630 6130
rect 48660 6050 48690 7160
rect 48730 7090 48790 7100
rect 48730 6120 48790 6130
rect 48820 6050 48850 7160
rect 48880 7090 48940 7100
rect 48880 6120 48940 6130
rect 48980 6050 49010 7160
rect 49040 7090 49100 7100
rect 49040 6120 49100 6130
rect 49130 6050 49160 7160
rect 49200 7090 49260 7100
rect 49200 6120 49260 6130
rect 49290 6050 49320 7160
rect 49360 7090 49420 7100
rect 49360 6120 49420 6130
rect 49450 6050 49480 7160
rect 49520 7090 49580 7100
rect 49520 6120 49580 6130
rect 49610 6050 49640 7160
rect 49670 7090 49730 7100
rect 49670 6120 49730 6130
rect 49760 6050 49790 7160
rect 49830 7090 49890 7100
rect 49830 6120 49890 6130
rect 49930 6050 49960 7160
rect 49990 7090 50050 7100
rect 49990 6120 50050 6130
rect 50080 6050 50110 7160
rect 50150 7090 50210 7100
rect 50150 6120 50210 6130
rect 50250 6050 50280 7160
rect 50350 7100 50520 7190
rect 50330 7090 50520 7100
rect 50330 6130 50340 7090
rect 50510 6800 50520 7090
rect 52520 6800 52920 8400
rect 71350 8310 71590 8700
rect 81910 8590 84010 8600
rect 81910 8350 81920 8590
rect 82300 8350 84010 8590
rect 81910 8340 84010 8350
rect 71190 8300 71870 8310
rect 71190 8100 71200 8300
rect 71860 8100 71870 8300
rect 71190 8090 71870 8100
rect 83660 8120 84010 8340
rect 66930 7960 73550 8050
rect 83660 7960 86150 8120
rect 66850 7900 66930 7910
rect 66850 6940 66860 7900
rect 66920 6940 66930 7900
rect 66850 6930 66930 6940
rect 66980 6860 67050 7960
rect 67110 7900 67190 7910
rect 67110 6940 67120 7900
rect 67180 6940 67190 7900
rect 67110 6930 67190 6940
rect 67240 6860 67310 7960
rect 67370 7900 67450 7910
rect 67370 6940 67380 7900
rect 67440 6940 67450 7900
rect 67370 6930 67450 6940
rect 67500 6860 67570 7960
rect 67630 7900 67710 7910
rect 67630 6940 67640 7900
rect 67700 6940 67710 7900
rect 67630 6930 67710 6940
rect 67760 6860 67830 7960
rect 67880 7900 67960 7910
rect 67880 6940 67890 7900
rect 67950 6940 67960 7900
rect 67880 6930 67960 6940
rect 50510 6400 52920 6800
rect 66930 6850 67110 6860
rect 67190 6850 67370 6860
rect 67450 6850 67630 6860
rect 67710 6850 67890 6860
rect 68010 6850 68080 7960
rect 68140 7900 68220 7910
rect 68140 6940 68150 7900
rect 68210 6940 68220 7900
rect 68140 6930 68220 6940
rect 68270 6850 68340 7960
rect 68400 7900 68480 7910
rect 68400 6940 68410 7900
rect 68470 6940 68480 7900
rect 68400 6930 68480 6940
rect 68530 6850 68600 7960
rect 68660 7900 68740 7910
rect 68660 6940 68670 7900
rect 68730 6940 68740 7900
rect 68660 6930 68740 6940
rect 68790 6850 68860 7960
rect 68910 7900 68990 7910
rect 68910 6940 68920 7900
rect 68980 6940 68990 7900
rect 68910 6930 68990 6940
rect 69050 6850 69120 7960
rect 69170 7900 69250 7910
rect 69170 6940 69180 7900
rect 69240 6940 69250 7900
rect 69170 6930 69250 6940
rect 69300 6850 69370 7960
rect 69430 7900 69510 7910
rect 69430 6940 69440 7900
rect 69500 6940 69510 7900
rect 69430 6930 69510 6940
rect 69560 6850 69630 7960
rect 69690 7900 69770 7910
rect 69690 6940 69700 7900
rect 69760 6940 69770 7900
rect 69690 6930 69770 6940
rect 69820 6850 69890 7960
rect 69950 7900 70030 7910
rect 69950 6940 69960 7900
rect 70020 7480 70030 7900
rect 70210 7900 70290 7910
rect 70210 7480 70220 7900
rect 70020 7340 70220 7480
rect 70020 6940 70030 7340
rect 69950 6930 70030 6940
rect 70210 6940 70220 7340
rect 70280 7480 70290 7900
rect 70450 7900 70530 7910
rect 70450 7480 70460 7900
rect 70280 7340 70460 7480
rect 70280 6940 70290 7340
rect 70210 6930 70290 6940
rect 70450 6940 70460 7340
rect 70520 6940 70530 7900
rect 70450 6930 70530 6940
rect 70590 6850 70660 7960
rect 70710 7900 70790 7910
rect 70710 6940 70720 7900
rect 70780 6940 70790 7900
rect 70710 6930 70790 6940
rect 70850 6850 70920 7960
rect 70970 7900 71050 7910
rect 70970 6940 70980 7900
rect 71040 6940 71050 7900
rect 70970 6930 71050 6940
rect 71100 6850 71170 7960
rect 71230 7900 71310 7910
rect 71230 6940 71240 7900
rect 71300 6940 71310 7900
rect 71230 6930 71310 6940
rect 71370 6850 71440 7960
rect 71490 7900 71570 7910
rect 71490 6940 71500 7900
rect 71560 6940 71570 7900
rect 71490 6930 71570 6940
rect 71620 6850 71690 7960
rect 71750 7900 71830 7910
rect 71750 6940 71760 7900
rect 71820 6940 71830 7900
rect 71750 6930 71830 6940
rect 71880 6850 71950 7960
rect 72000 7900 72080 7910
rect 72000 6940 72010 7900
rect 72070 6940 72080 7900
rect 72000 6930 72080 6940
rect 72140 6850 72210 7960
rect 72260 7900 72340 7910
rect 72260 6940 72270 7900
rect 72330 6940 72340 7900
rect 72260 6930 72340 6940
rect 72400 6850 72470 7960
rect 72520 7900 72600 7910
rect 72520 6940 72530 7900
rect 72590 6940 72600 7900
rect 72520 6930 72600 6940
rect 72660 6850 72730 7960
rect 72780 7900 72860 7910
rect 72780 6940 72790 7900
rect 72850 6940 72860 7900
rect 72780 6930 72860 6940
rect 72920 6850 72990 7960
rect 73040 7900 73120 7910
rect 73040 6940 73050 7900
rect 73110 6940 73120 7900
rect 73040 6930 73120 6940
rect 73170 6850 73240 7960
rect 73300 7900 73380 7910
rect 73300 6940 73310 7900
rect 73370 6940 73380 7900
rect 73300 6930 73380 6940
rect 73430 6850 73500 7960
rect 73560 7900 73640 7910
rect 73560 6940 73570 7900
rect 73630 6940 73640 7900
rect 73560 6930 73640 6940
rect 66930 6720 73550 6850
rect 83660 6780 84010 7960
rect 84290 7900 86150 7960
rect 84250 7820 84310 7830
rect 84250 6860 84310 6870
rect 84400 7820 84460 7830
rect 84400 6860 84460 6870
rect 84560 7820 84620 7830
rect 84560 6860 84620 6870
rect 84720 7820 84780 7830
rect 84720 6860 84780 6870
rect 84880 7820 84940 7830
rect 84880 6860 84940 6870
rect 85030 7820 85090 7830
rect 85030 6860 85090 6870
rect 85190 7820 85250 7830
rect 85190 6860 85250 6870
rect 85350 7820 85410 7830
rect 85350 6860 85410 6870
rect 85510 7820 85570 7830
rect 85510 6860 85570 6870
rect 85670 7820 85730 7830
rect 85670 6860 85730 6870
rect 85820 7820 85880 7830
rect 85820 6860 85880 6870
rect 85980 7820 86040 7830
rect 85980 6860 86040 6870
rect 86140 7820 86200 7830
rect 86140 6860 86200 6870
rect 50510 6130 50520 6400
rect 50330 6120 50520 6130
rect 48180 6000 48230 6050
rect 48330 6000 48380 6050
rect 48810 6000 48860 6050
rect 48970 6000 49020 6050
rect 49440 6000 49490 6050
rect 49600 6000 49650 6050
rect 50070 6000 50120 6050
rect 50240 6000 50290 6050
rect 50350 6030 50520 6120
rect 52520 6330 52920 6400
rect 66850 6660 66930 6670
rect 52520 6320 53300 6330
rect 47840 5990 51280 6000
rect 47840 5810 50720 5990
rect 51270 5810 51280 5990
rect 52520 5920 52530 6320
rect 53290 5920 53300 6320
rect 52520 5910 53300 5920
rect 47840 5800 51280 5810
rect 66850 5700 66860 6660
rect 66920 5700 66930 6660
rect 66850 5690 66930 5700
rect 66980 5620 67050 6720
rect 67110 6660 67190 6670
rect 67110 5700 67120 6660
rect 67180 5700 67190 6660
rect 67110 5690 67190 5700
rect 67240 5620 67310 6720
rect 67370 6660 67450 6670
rect 67370 5700 67380 6660
rect 67440 5700 67450 6660
rect 67370 5690 67450 5700
rect 67500 5620 67570 6720
rect 67630 6660 67710 6670
rect 67630 5700 67640 6660
rect 67700 5700 67710 6660
rect 67630 5690 67710 5700
rect 67760 5620 67830 6720
rect 67880 6660 67960 6670
rect 67880 5700 67890 6660
rect 67950 5700 67960 6660
rect 67880 5690 67960 5700
rect 68010 5620 68080 6720
rect 68140 6660 68220 6670
rect 68140 5700 68150 6660
rect 68210 5700 68220 6660
rect 68140 5690 68220 5700
rect 68270 5620 68340 6720
rect 68400 6660 68480 6670
rect 68400 5700 68410 6660
rect 68470 5700 68480 6660
rect 68400 5690 68480 5700
rect 68530 5620 68600 6720
rect 68660 6660 68740 6670
rect 68660 5700 68670 6660
rect 68730 5700 68740 6660
rect 68660 5690 68740 5700
rect 68790 5620 68860 6720
rect 68910 6660 68990 6670
rect 68910 5700 68920 6660
rect 68980 5700 68990 6660
rect 68910 5690 68990 5700
rect 69050 5620 69120 6720
rect 69170 6660 69250 6670
rect 69170 5700 69180 6660
rect 69240 5700 69250 6660
rect 69170 5690 69250 5700
rect 69300 5620 69370 6720
rect 69430 6660 69510 6670
rect 69430 5700 69440 6660
rect 69500 5700 69510 6660
rect 69430 5690 69510 5700
rect 69560 5620 69630 6720
rect 69690 6660 69770 6670
rect 69690 5700 69700 6660
rect 69760 5700 69770 6660
rect 69690 5690 69770 5700
rect 69820 5620 69890 6720
rect 69950 6660 70030 6670
rect 69950 5700 69960 6660
rect 70020 5700 70030 6660
rect 69950 5690 70030 5700
rect 70080 6660 70400 6720
rect 70080 5700 70220 6660
rect 70280 5700 70400 6660
rect 70080 5620 70400 5700
rect 70450 6660 70530 6670
rect 70450 5700 70460 6660
rect 70520 5700 70530 6660
rect 70450 5690 70530 5700
rect 70590 5620 70660 6720
rect 70710 6660 70790 6670
rect 70710 5700 70720 6660
rect 70780 5700 70790 6660
rect 70710 5690 70790 5700
rect 70850 5620 70920 6720
rect 70970 6660 71050 6670
rect 70970 5700 70980 6660
rect 71040 5700 71050 6660
rect 70970 5690 71050 5700
rect 71100 5620 71170 6720
rect 71230 6660 71310 6670
rect 71230 5700 71240 6660
rect 71300 5700 71310 6660
rect 71230 5690 71310 5700
rect 71370 5620 71440 6720
rect 71490 6660 71570 6670
rect 71490 5700 71500 6660
rect 71560 5700 71570 6660
rect 71490 5690 71570 5700
rect 71620 5620 71690 6720
rect 71750 6660 71830 6670
rect 71750 5700 71760 6660
rect 71820 5700 71830 6660
rect 71750 5690 71830 5700
rect 71880 5620 71950 6720
rect 72000 6660 72080 6670
rect 72000 5700 72010 6660
rect 72070 5700 72080 6660
rect 72000 5690 72080 5700
rect 72140 5620 72210 6720
rect 72260 6660 72340 6670
rect 72260 5700 72270 6660
rect 72330 5700 72340 6660
rect 72260 5690 72340 5700
rect 72400 5620 72470 6720
rect 72520 6660 72600 6670
rect 72520 5700 72530 6660
rect 72590 5700 72600 6660
rect 72520 5690 72600 5700
rect 72660 5620 72730 6720
rect 72780 6660 72860 6670
rect 72780 5700 72790 6660
rect 72850 5700 72860 6660
rect 72780 5690 72860 5700
rect 72920 5620 72990 6720
rect 73040 6660 73120 6670
rect 73040 5700 73050 6660
rect 73110 5700 73120 6660
rect 73040 5690 73120 5700
rect 73170 5620 73240 6720
rect 73300 6660 73380 6670
rect 73300 5700 73310 6660
rect 73370 5700 73380 6660
rect 73300 5690 73380 5700
rect 73430 5620 73500 6720
rect 83660 6670 83770 6780
rect 84000 6670 84010 6780
rect 73560 6660 73640 6670
rect 73560 5700 73570 6660
rect 73630 5700 73640 6660
rect 73560 5690 73640 5700
rect 66930 5490 73550 5620
rect 83660 5490 84010 6670
rect 84310 6780 86140 6790
rect 84310 6670 84670 6780
rect 84830 6670 86140 6780
rect 84310 6660 86140 6670
rect 84250 6580 84310 6590
rect 84250 5620 84310 5630
rect 84400 6580 84460 6590
rect 84400 5620 84460 5630
rect 84560 6580 84620 6590
rect 84560 5620 84620 5630
rect 84720 6580 84780 6590
rect 84720 5620 84780 5630
rect 84880 6580 84940 6590
rect 84880 5620 84940 5630
rect 85030 6580 85090 6590
rect 85030 5620 85090 5630
rect 85190 6580 85250 6590
rect 85190 5620 85250 5630
rect 85350 6580 85410 6590
rect 85350 5620 85410 5630
rect 85510 6580 85570 6590
rect 85510 5620 85570 5630
rect 85670 6580 85730 6590
rect 85670 5620 85730 5630
rect 85820 6580 85880 6590
rect 85820 5620 85880 5630
rect 85980 6580 86040 6590
rect 85980 5620 86040 5630
rect 86140 6580 86200 6590
rect 86140 5620 86200 5630
rect 84270 5490 86150 5560
rect 13960 5120 14260 5130
rect 47480 5280 47800 5290
rect 13960 4820 14100 5120
rect 47480 5100 47490 5280
rect 47790 5100 47800 5280
rect 47480 5090 47800 5100
rect 66850 5420 66930 5430
rect 8720 4740 10080 4820
rect 12780 4740 14100 4820
rect 47740 4460 51240 4600
rect 39080 4310 45720 4450
rect 47740 4430 51010 4460
rect 38770 3700 39070 4270
rect 38770 3690 39090 3700
rect 38830 3310 39030 3690
rect 38770 3300 39090 3310
rect 38770 3040 39000 3300
rect 39150 3240 39230 4310
rect 39280 4250 39360 4260
rect 39280 3310 39290 4250
rect 39350 3310 39360 4250
rect 39280 3300 39360 3310
rect 39410 3240 39490 4310
rect 39540 3690 39600 3700
rect 39540 3300 39600 3310
rect 39660 3240 39740 4310
rect 39790 4250 39870 4260
rect 39790 3310 39800 4250
rect 39860 3310 39870 4250
rect 39790 3300 39870 3310
rect 39920 3240 40000 4310
rect 40060 3690 40120 3700
rect 40060 3300 40120 3310
rect 40180 3240 40260 4310
rect 40310 4240 40390 4260
rect 40310 3310 40320 4240
rect 40380 3310 40390 4240
rect 40310 3300 40390 3310
rect 40430 3240 40510 4310
rect 40580 3690 40640 3700
rect 40580 3300 40640 3310
rect 40700 3240 40780 4310
rect 40820 4250 40900 4260
rect 40820 3310 40830 4250
rect 40890 3310 40900 4250
rect 40820 3300 40900 3310
rect 40950 3240 41030 4310
rect 41090 3690 41150 3700
rect 41090 3300 41150 3310
rect 41210 3240 41290 4310
rect 41340 4250 41420 4260
rect 41340 3310 41350 4250
rect 41410 3310 41420 4250
rect 41340 3300 41420 3310
rect 41470 3240 41550 4310
rect 41610 3690 41670 3700
rect 41610 3300 41670 3310
rect 41730 3240 41810 4310
rect 41860 4250 41940 4260
rect 41860 3310 41870 4250
rect 41930 3310 41940 4250
rect 41860 3300 41940 3310
rect 41990 3240 42070 4310
rect 42120 3690 42180 3700
rect 42120 3300 42180 3310
rect 42250 3240 42330 4310
rect 42370 4250 42450 4260
rect 42370 3310 42380 4250
rect 42440 3310 42450 4250
rect 42370 3300 42450 3310
rect 42500 3240 42580 4310
rect 42640 3690 42700 3700
rect 42640 3300 42700 3310
rect 42760 3240 42840 4310
rect 42890 4250 42970 4260
rect 42890 3310 42900 4250
rect 42960 3310 42970 4250
rect 42890 3300 42970 3310
rect 43020 3240 43100 4310
rect 43160 3690 43220 3700
rect 43160 3300 43220 3310
rect 43280 3240 43360 4310
rect 43400 4250 43480 4260
rect 43400 3310 43410 4250
rect 43470 3310 43480 4250
rect 43400 3300 43480 3310
rect 43540 3240 43620 4310
rect 43670 3690 43730 3700
rect 43670 3300 43730 3310
rect 43790 3240 43870 4310
rect 43920 4250 44000 4260
rect 43920 3310 43930 4250
rect 43990 3310 44000 4250
rect 43920 3300 44000 3310
rect 44050 3240 44130 4310
rect 44190 3690 44250 3700
rect 44190 3300 44250 3310
rect 44310 3240 44390 4310
rect 44440 4250 44520 4260
rect 44440 3310 44450 4250
rect 44510 3310 44520 4250
rect 44440 3300 44520 3310
rect 44570 3240 44650 4310
rect 44700 3690 44760 3700
rect 44700 3300 44760 3310
rect 44820 3240 44900 4310
rect 44950 4250 45030 4260
rect 44950 3310 44960 4250
rect 45020 3310 45030 4250
rect 44950 3300 45030 3310
rect 45080 3240 45160 4310
rect 45220 3690 45280 3700
rect 45220 3300 45280 3310
rect 45340 3240 45420 4310
rect 45470 4250 45550 4260
rect 45470 3310 45480 4250
rect 45540 3310 45550 4250
rect 45470 3300 45550 3310
rect 45600 3240 45680 4310
rect 45750 3700 46040 4270
rect 47140 4210 47220 4220
rect 45740 3690 46050 3700
rect 45800 3310 45990 3690
rect 45740 3300 45800 3310
rect 45830 3300 46050 3310
rect 39090 3230 45740 3240
rect 39090 3110 39100 3230
rect 39240 3110 39400 3230
rect 39750 3110 39910 3230
rect 40260 3110 40430 3230
rect 40780 3110 40940 3230
rect 41290 3110 41460 3230
rect 41810 3110 41980 3230
rect 42330 3110 42490 3230
rect 42840 3110 43010 3230
rect 43360 3110 43520 3230
rect 43870 3110 44040 3230
rect 44390 3110 44560 3230
rect 44910 3110 45070 3230
rect 45420 3110 45590 3230
rect 45730 3110 45740 3230
rect 39090 3100 45740 3110
rect 38770 2480 39080 3040
rect 38770 2470 39090 2480
rect 38830 2090 39030 2470
rect 38770 2080 39090 2090
rect 39150 2020 39230 3100
rect 39280 3030 39360 3040
rect 39280 2090 39290 3030
rect 39350 2090 39360 3030
rect 39280 2080 39360 2090
rect 39410 2020 39490 3100
rect 39540 2470 39600 2480
rect 39540 2080 39600 2090
rect 39660 2020 39740 3100
rect 39790 3030 39870 3040
rect 39790 2090 39800 3030
rect 39860 2090 39870 3030
rect 39790 2080 39870 2090
rect 39920 2020 40000 3100
rect 40060 2470 40120 2480
rect 40060 2080 40120 2090
rect 40180 2020 40260 3100
rect 40310 3030 40390 3040
rect 40310 2090 40320 3030
rect 40380 2090 40390 3030
rect 40310 2080 40390 2090
rect 40430 2020 40510 3100
rect 40580 2470 40640 2480
rect 40580 2080 40640 2090
rect 40700 2020 40780 3100
rect 40820 3030 40900 3040
rect 40820 2090 40830 3030
rect 40890 2090 40900 3030
rect 40820 2080 40900 2090
rect 40950 2020 41030 3100
rect 41090 2470 41150 2480
rect 41090 2080 41150 2090
rect 41210 2020 41550 3100
rect 41610 2470 41670 2480
rect 41610 2080 41670 2090
rect 41730 2020 41810 3100
rect 41860 3030 41940 3040
rect 41860 2090 41870 3030
rect 41930 2090 41940 3030
rect 41860 2080 41940 2090
rect 41990 2020 42070 3100
rect 42120 2470 42180 2480
rect 42120 2080 42180 2090
rect 42250 2020 42330 3100
rect 42370 3030 42450 3040
rect 42370 2090 42380 3030
rect 42440 2090 42450 3030
rect 42370 2080 42450 2090
rect 42500 2020 42580 3100
rect 42640 2470 42700 2480
rect 42640 2080 42700 2090
rect 42760 2020 42840 3100
rect 42890 3030 42970 3040
rect 42890 2090 42900 3030
rect 42960 2090 42970 3030
rect 42890 2080 42970 2090
rect 43020 2020 43100 3100
rect 43160 2470 43220 2480
rect 43160 2080 43220 2090
rect 43280 2020 43360 3100
rect 43400 3030 43480 3040
rect 43400 2090 43410 3030
rect 43470 2090 43480 3030
rect 43400 2080 43480 2090
rect 43540 2020 43620 3100
rect 43670 2470 43730 2480
rect 43670 2080 43730 2090
rect 43790 2020 43870 3100
rect 43920 3030 44000 3040
rect 43920 2090 43930 3030
rect 43990 2090 44000 3030
rect 43920 2080 44000 2090
rect 44050 2020 44130 3100
rect 44190 2470 44250 2480
rect 44190 2080 44250 2090
rect 44310 2020 44390 3100
rect 44440 3030 44520 3040
rect 44440 2090 44450 3030
rect 44510 2090 44520 3030
rect 44440 2080 44520 2090
rect 44570 2020 44650 3100
rect 44700 2470 44760 2480
rect 44700 2080 44760 2090
rect 44820 2020 44900 3100
rect 44950 3030 45030 3040
rect 44950 2090 44960 3030
rect 45020 2090 45030 3030
rect 44950 2080 45030 2090
rect 45080 2020 45160 3100
rect 45220 2470 45280 2480
rect 45220 2080 45280 2090
rect 45340 2020 45420 3100
rect 45470 3030 45550 3040
rect 45470 2090 45480 3030
rect 45540 2090 45550 3030
rect 45470 2080 45550 2090
rect 45600 2020 45680 3100
rect 45830 3040 46040 3300
rect 47140 3250 47150 4210
rect 47210 3250 47220 4210
rect 47140 3240 47220 3250
rect 47270 4210 47620 4310
rect 47740 4280 48180 4430
rect 47270 3250 47420 4210
rect 47480 3250 47620 4210
rect 45750 2480 46040 3040
rect 47140 2980 47220 2990
rect 45740 2470 46050 2480
rect 45800 2090 45990 2470
rect 45740 2080 46050 2090
rect 47140 2020 47150 2980
rect 47210 2020 47220 2980
rect 39090 1940 45730 2020
rect 47140 2010 47220 2020
rect 47270 2980 47620 3250
rect 47660 4210 47740 4220
rect 47660 3250 47670 4210
rect 47730 3250 47740 4210
rect 47660 3240 47740 3250
rect 47270 2020 47420 2980
rect 47480 2020 47620 2980
rect 39090 1880 45740 1940
rect 47270 1920 47620 2020
rect 47660 2980 47740 2990
rect 47660 2020 47670 2980
rect 47730 2020 47740 2980
rect 47660 2010 47740 2020
rect 47790 1920 47880 4280
rect 47920 4210 48000 4220
rect 47920 3250 47930 4210
rect 47990 3250 48000 4210
rect 47920 3240 48000 3250
rect 47920 2980 48000 2990
rect 47920 2020 47930 2980
rect 47990 2020 48000 2980
rect 47920 2010 48000 2020
rect 48040 1920 48130 4280
rect 48180 4210 48260 4220
rect 48180 3250 48190 4210
rect 48250 3250 48260 4210
rect 48180 3240 48260 3250
rect 48300 4210 48650 4310
rect 48780 4280 49220 4430
rect 48300 3250 48450 4210
rect 48510 3250 48650 4210
rect 48180 2980 48260 2990
rect 48180 2020 48190 2980
rect 48250 2020 48260 2980
rect 48180 2010 48260 2020
rect 48300 2980 48650 3250
rect 48690 4210 48770 4220
rect 48690 3250 48700 4210
rect 48760 3250 48770 4210
rect 48690 3240 48770 3250
rect 48300 2020 48450 2980
rect 48510 2020 48650 2980
rect 48300 1920 48650 2020
rect 48690 2980 48770 2990
rect 48690 2020 48700 2980
rect 48760 2020 48770 2980
rect 48690 2010 48770 2020
rect 48820 1920 48910 4280
rect 48950 4210 49030 4220
rect 48950 3250 48960 4210
rect 49020 3250 49030 4210
rect 48950 3240 49030 3250
rect 48950 2980 49030 2990
rect 48950 2020 48960 2980
rect 49020 2020 49030 2980
rect 48950 2010 49030 2020
rect 49080 1920 49170 4280
rect 49210 4210 49290 4220
rect 49210 3250 49220 4210
rect 49280 3250 49290 4210
rect 49210 3240 49290 3250
rect 49330 4210 49680 4310
rect 49800 4280 50240 4430
rect 49330 3250 49480 4210
rect 49540 3250 49680 4210
rect 49210 2980 49290 2990
rect 49210 2020 49220 2980
rect 49280 2020 49290 2980
rect 49210 2010 49290 2020
rect 49330 2980 49680 3250
rect 49730 4210 49810 4220
rect 49730 3250 49740 4210
rect 49800 3250 49810 4210
rect 49730 3240 49810 3250
rect 49330 2020 49480 2980
rect 49540 2020 49680 2980
rect 49330 1920 49680 2020
rect 49730 2980 49810 2990
rect 49730 2020 49740 2980
rect 49800 2020 49810 2980
rect 49730 2010 49810 2020
rect 49850 1920 49940 4280
rect 49980 4210 50060 4220
rect 49980 3250 49990 4210
rect 50050 3250 50060 4210
rect 49980 3240 50060 3250
rect 49980 2980 50060 2990
rect 49980 2020 49990 2980
rect 50050 2020 50060 2980
rect 49980 2010 50060 2020
rect 50110 1920 50200 4280
rect 50250 4210 50330 4220
rect 50250 3250 50260 4210
rect 50320 3250 50330 4210
rect 51000 4070 51010 4430
rect 51230 4070 51240 4460
rect 66850 4460 66860 5420
rect 66920 4460 66930 5420
rect 66850 4450 66930 4460
rect 66980 4380 67050 5490
rect 67110 5420 67190 5430
rect 67110 4460 67120 5420
rect 67180 4460 67190 5420
rect 67110 4450 67190 4460
rect 67240 4380 67310 5490
rect 67370 5420 67450 5430
rect 67370 4460 67380 5420
rect 67440 4460 67450 5420
rect 67370 4450 67450 4460
rect 67500 4380 67570 5490
rect 67630 5420 67710 5430
rect 67630 4460 67640 5420
rect 67700 4460 67710 5420
rect 67630 4450 67710 4460
rect 67760 4380 67830 5490
rect 67880 5420 67960 5430
rect 67880 4460 67890 5420
rect 67950 4460 67960 5420
rect 67880 4450 67960 4460
rect 68010 4380 68080 5490
rect 68140 5420 68220 5430
rect 68140 4460 68150 5420
rect 68210 4460 68220 5420
rect 68140 4450 68220 4460
rect 68270 4380 68340 5490
rect 68400 5420 68480 5430
rect 68400 4460 68410 5420
rect 68470 4460 68480 5420
rect 68400 4450 68480 4460
rect 68530 4380 68600 5490
rect 68660 5420 68740 5430
rect 68660 4460 68670 5420
rect 68730 4460 68740 5420
rect 68660 4450 68740 4460
rect 68790 4380 68860 5490
rect 68910 5420 68990 5430
rect 68910 4460 68920 5420
rect 68980 4460 68990 5420
rect 68910 4450 68990 4460
rect 69050 4380 69120 5490
rect 69170 5420 69250 5430
rect 69170 4460 69180 5420
rect 69240 4460 69250 5420
rect 69170 4450 69250 4460
rect 69300 4380 69370 5490
rect 69430 5420 69510 5430
rect 69430 4460 69440 5420
rect 69500 4460 69510 5420
rect 69430 4450 69510 4460
rect 69560 4380 69630 5490
rect 69690 5420 69770 5430
rect 69690 4460 69700 5420
rect 69760 4460 69770 5420
rect 69690 4450 69770 4460
rect 69820 4380 69890 5490
rect 69950 5420 70030 5430
rect 69950 4460 69960 5420
rect 70020 4460 70030 5420
rect 69950 4450 70030 4460
rect 70080 5420 70400 5490
rect 70080 4460 70220 5420
rect 70280 4460 70400 5420
rect 70080 4380 70400 4460
rect 70450 5420 70530 5430
rect 70450 4460 70460 5420
rect 70520 4460 70530 5420
rect 70450 4450 70530 4460
rect 70590 4380 70660 5490
rect 70710 5420 70790 5430
rect 70710 4460 70720 5420
rect 70780 4460 70790 5420
rect 70710 4450 70790 4460
rect 70850 4380 70920 5490
rect 70970 5420 71050 5430
rect 70970 4460 70980 5420
rect 71040 4460 71050 5420
rect 70970 4450 71050 4460
rect 71100 4380 71170 5490
rect 71230 5420 71310 5430
rect 71230 4460 71240 5420
rect 71300 4460 71310 5420
rect 71230 4450 71310 4460
rect 71370 4380 71440 5490
rect 71490 5420 71570 5430
rect 71490 4460 71500 5420
rect 71560 4460 71570 5420
rect 71490 4450 71570 4460
rect 71620 4380 71690 5490
rect 71750 5420 71830 5430
rect 71750 4460 71760 5420
rect 71820 4460 71830 5420
rect 71750 4450 71830 4460
rect 71880 4380 71950 5490
rect 72000 5420 72080 5430
rect 72000 4460 72010 5420
rect 72070 4460 72080 5420
rect 72000 4450 72080 4460
rect 72140 4380 72210 5490
rect 72260 5420 72340 5430
rect 72260 4460 72270 5420
rect 72330 4460 72340 5420
rect 72260 4450 72340 4460
rect 72400 4380 72470 5490
rect 72520 5420 72600 5430
rect 72520 4460 72530 5420
rect 72590 4460 72600 5420
rect 72520 4450 72600 4460
rect 72660 4380 72730 5490
rect 72780 5420 72860 5430
rect 72780 4460 72790 5420
rect 72850 4460 72860 5420
rect 72780 4450 72860 4460
rect 72920 4380 72990 5490
rect 73040 5420 73120 5430
rect 73040 4460 73050 5420
rect 73110 4460 73120 5420
rect 73040 4450 73120 4460
rect 73170 4380 73240 5490
rect 73300 5420 73380 5430
rect 73300 4460 73310 5420
rect 73370 4460 73380 5420
rect 73300 4450 73380 4460
rect 73430 4380 73500 5490
rect 73560 5420 73640 5430
rect 73560 4460 73570 5420
rect 73630 4460 73640 5420
rect 83660 5370 86150 5490
rect 84320 4650 86610 4780
rect 84320 4570 86130 4650
rect 73560 4450 73640 4460
rect 84240 4490 84300 4500
rect 66930 4250 73550 4380
rect 51000 4060 51240 4070
rect 66850 4180 66930 4190
rect 50250 3240 50330 3250
rect 66850 3220 66860 4180
rect 66920 3220 66930 4180
rect 66850 3210 66930 3220
rect 66980 3140 67050 4250
rect 67110 4180 67190 4190
rect 67110 3220 67120 4180
rect 67180 3220 67190 4180
rect 67110 3210 67190 3220
rect 67240 3140 67310 4250
rect 67370 4180 67450 4190
rect 67370 3220 67380 4180
rect 67440 3220 67450 4180
rect 67370 3210 67450 3220
rect 67500 3140 67570 4250
rect 67630 4180 67710 4190
rect 67630 3220 67640 4180
rect 67700 3220 67710 4180
rect 67630 3210 67710 3220
rect 67760 3140 67830 4250
rect 67880 4180 67960 4190
rect 67880 3220 67890 4180
rect 67950 3220 67960 4180
rect 67880 3210 67960 3220
rect 68010 3140 68080 4250
rect 68140 4180 68220 4190
rect 68140 3220 68150 4180
rect 68210 3220 68220 4180
rect 68140 3210 68220 3220
rect 68270 3140 68340 4250
rect 68400 4180 68480 4190
rect 68400 3220 68410 4180
rect 68470 3220 68480 4180
rect 68400 3210 68480 3220
rect 68530 3140 68600 4250
rect 68660 4180 68740 4190
rect 68660 3220 68670 4180
rect 68730 3220 68740 4180
rect 68660 3210 68740 3220
rect 68790 3140 68860 4250
rect 68910 4180 68990 4190
rect 68910 3220 68920 4180
rect 68980 3220 68990 4180
rect 68910 3210 68990 3220
rect 69050 3140 69120 4250
rect 69170 4180 69250 4190
rect 69170 3220 69180 4180
rect 69240 3220 69250 4180
rect 69170 3210 69250 3220
rect 69300 3140 69370 4250
rect 69430 4180 69510 4190
rect 69430 3220 69440 4180
rect 69500 3220 69510 4180
rect 69430 3210 69510 3220
rect 69560 3140 69630 4250
rect 69690 4180 69770 4190
rect 69690 3220 69700 4180
rect 69760 3220 69770 4180
rect 69690 3210 69770 3220
rect 69820 3140 69890 4250
rect 69950 4180 70030 4190
rect 69950 3220 69960 4180
rect 70020 3220 70030 4180
rect 69950 3210 70030 3220
rect 70080 4180 70400 4250
rect 70080 3220 70220 4180
rect 70280 3220 70400 4180
rect 70080 3140 70400 3220
rect 70450 4180 70530 4190
rect 70450 3220 70460 4180
rect 70520 3220 70530 4180
rect 70450 3210 70530 3220
rect 70590 3140 70660 4250
rect 70710 4180 70790 4190
rect 70710 3220 70720 4180
rect 70780 3220 70790 4180
rect 70710 3210 70790 3220
rect 70850 3140 70920 4250
rect 70970 4180 71050 4190
rect 70970 3220 70980 4180
rect 71040 3220 71050 4180
rect 70970 3210 71050 3220
rect 71100 3140 71170 4250
rect 71230 4180 71310 4190
rect 71230 3220 71240 4180
rect 71300 3220 71310 4180
rect 71230 3210 71310 3220
rect 71370 3140 71440 4250
rect 71490 4180 71570 4190
rect 71490 3220 71500 4180
rect 71560 3220 71570 4180
rect 71490 3210 71570 3220
rect 71620 3140 71690 4250
rect 71750 4180 71830 4190
rect 71750 3220 71760 4180
rect 71820 3220 71830 4180
rect 71750 3210 71830 3220
rect 71880 3140 71950 4250
rect 72000 4180 72080 4190
rect 72000 3220 72010 4180
rect 72070 3220 72080 4180
rect 72000 3210 72080 3220
rect 72140 3140 72210 4250
rect 72260 4180 72340 4190
rect 72260 3220 72270 4180
rect 72330 3220 72340 4180
rect 72260 3210 72340 3220
rect 72400 3140 72470 4250
rect 72520 4180 72600 4190
rect 72520 3220 72530 4180
rect 72590 3220 72600 4180
rect 72520 3210 72600 3220
rect 72660 3140 72730 4250
rect 72780 4180 72860 4190
rect 72780 3220 72790 4180
rect 72850 3220 72860 4180
rect 72780 3210 72860 3220
rect 72920 3140 72990 4250
rect 73040 4180 73120 4190
rect 73040 3220 73050 4180
rect 73110 3220 73120 4180
rect 73040 3210 73120 3220
rect 73170 3140 73240 4250
rect 73300 4180 73380 4190
rect 73300 3220 73310 4180
rect 73370 3220 73380 4180
rect 73300 3210 73380 3220
rect 73430 3140 73500 4250
rect 73560 4180 73640 4190
rect 73560 3220 73570 4180
rect 73630 3220 73640 4180
rect 84240 3530 84300 3540
rect 84390 4490 84450 4500
rect 84390 3530 84450 3540
rect 84550 4490 84610 4500
rect 84550 3530 84610 3540
rect 84710 4490 84770 4500
rect 84710 3530 84770 3540
rect 84870 4490 84930 4500
rect 84870 3530 84930 3540
rect 85020 4490 85080 4500
rect 85020 3530 85080 3540
rect 85180 4490 85240 4500
rect 85180 3530 85240 3540
rect 85340 4490 85400 4500
rect 85340 3530 85400 3540
rect 85500 4490 85560 4500
rect 85500 3530 85560 3540
rect 85660 4490 85720 4500
rect 85660 3530 85720 3540
rect 85810 4490 85870 4500
rect 85810 3530 85870 3540
rect 85970 4490 86030 4500
rect 85970 3530 86030 3540
rect 86130 4490 86190 4500
rect 86130 3530 86190 3540
rect 84300 3340 86110 3470
rect 86400 3270 86610 4650
rect 73560 3210 73640 3220
rect 84240 3260 84300 3270
rect 66930 3070 73550 3140
rect 50250 2980 50330 2990
rect 50250 2020 50260 2980
rect 50320 2020 50330 2980
rect 84240 2300 84300 2310
rect 84390 3260 84450 3270
rect 84390 2300 84450 2310
rect 84550 3260 84610 3270
rect 84550 2300 84610 2310
rect 84710 3260 84770 3270
rect 84710 2300 84770 2310
rect 84870 3260 84930 3270
rect 84870 2300 84930 2310
rect 85020 3260 85080 3270
rect 85020 2300 85080 2310
rect 85180 3260 85240 3270
rect 85180 2300 85240 2310
rect 85340 3260 85400 3270
rect 85340 2300 85400 2310
rect 85500 3260 85560 3270
rect 85500 2300 85560 2310
rect 85660 3260 85720 3270
rect 85660 2300 85720 2310
rect 85810 3260 85870 3270
rect 85810 2300 85870 2310
rect 85970 3260 86030 3270
rect 85970 2300 86030 2310
rect 86130 3260 86190 3270
rect 86130 2300 86190 2310
rect 86400 3260 93630 3270
rect 86400 2870 93240 3260
rect 93620 2870 93630 3260
rect 86400 2860 93630 2870
rect 84310 2160 86110 2230
rect 86400 2160 86610 2860
rect 84310 2020 86610 2160
rect 50250 2010 50330 2020
rect 39100 1560 39260 1880
rect 39560 1560 39720 1880
rect 40080 1560 40240 1880
rect 40600 1560 40760 1880
rect 41060 1560 41220 1880
rect 41560 1560 41720 1880
rect 42040 1560 42200 1880
rect 42560 1560 42720 1880
rect 43000 1560 43160 1880
rect 43580 1560 43740 1880
rect 44140 1560 44300 1880
rect 44580 1560 44740 1880
rect 44980 1560 45140 1880
rect 45580 1560 45740 1880
rect 7780 1480 45740 1560
rect 7770 920 45740 1480
rect 51540 1080 52570 1140
rect 51540 930 51610 1080
rect 51350 920 51610 930
rect 7770 400 8320 920
rect 51350 710 51360 920
rect 51590 780 51610 920
rect 51780 1010 52050 1020
rect 52510 1010 52570 1080
rect 53390 1030 53630 1040
rect 51780 850 51790 1010
rect 52040 850 52050 1010
rect 53390 970 53400 1030
rect 52110 960 52510 970
rect 52110 900 52190 960
rect 52420 900 52510 960
rect 52110 890 52510 900
rect 52580 960 53400 970
rect 52580 900 52680 960
rect 52830 900 53400 960
rect 52580 890 53400 900
rect 51780 840 52050 850
rect 52510 780 52570 850
rect 53390 840 53400 890
rect 53620 840 53630 1030
rect 53390 830 53630 840
rect 51590 710 52570 780
rect 51350 700 52570 710
rect 7180 390 8780 400
rect 7180 10 7190 390
rect 8770 10 8780 390
rect 7180 0 8780 10
<< via1 >>
rect 3000 44840 3080 45140
rect 3550 44840 3630 45140
rect 4110 44840 4190 45140
rect 4660 44840 4740 45140
rect 5210 44840 5290 45140
rect 5770 44840 5850 45140
rect 6320 44840 6400 45140
rect 6870 44840 6950 45140
rect 7410 44840 7490 45140
rect 7970 44840 8050 45140
rect 8510 44840 8590 45140
rect 9070 44840 9150 45140
rect 9620 44840 9700 45140
rect 10180 44840 10260 45140
rect 10730 44840 10810 45140
rect 11290 44840 11370 45140
rect 11890 44770 12140 44960
rect 12390 44840 12470 45140
rect 12940 44840 13020 45140
rect 13480 44840 13560 45140
rect 14040 44840 14120 45140
rect 14590 44840 14670 45140
rect 15140 44840 15220 45140
rect 16250 44840 16330 45140
rect 16800 44840 16880 45140
rect 17350 44840 17430 45140
rect 17910 44840 17990 45140
rect 18460 44840 18540 45140
rect 19010 44840 19090 45140
rect 19560 44840 19640 45140
rect 20120 44840 20200 45140
rect 20670 44840 20750 45140
rect 21220 44840 21300 45140
rect 21770 44840 21850 45140
rect 22310 44840 22390 45140
rect 23980 44840 24060 45140
rect 24480 44960 24650 45140
rect 3510 44440 3640 44580
rect 25580 44960 25750 45140
rect 27010 44870 27210 45010
rect 28110 44450 28360 44620
rect 70610 12770 70980 12960
rect 66330 12500 66560 12690
rect 66960 12500 67190 12690
rect 66250 11450 66310 12420
rect 66250 10210 66310 11180
rect 66420 11450 66480 12420
rect 66420 10210 66480 11180
rect 66570 11450 66630 12420
rect 66570 10210 66630 11180
rect 66730 11450 66790 12420
rect 66730 10210 66790 11180
rect 66890 11450 66950 12420
rect 66890 10210 66950 11180
rect 67050 11450 67110 12420
rect 67050 10210 67110 11180
rect 67600 12500 67830 12690
rect 67200 11450 67260 12420
rect 67200 10210 67260 11180
rect 53010 9490 53280 10090
rect 66650 9940 66870 10130
rect 67360 11450 67420 12420
rect 67360 10210 67420 11180
rect 67520 11450 67580 12420
rect 67520 10210 67580 11180
rect 67680 11450 67740 12420
rect 67680 10210 67740 11180
rect 68230 12500 68460 12690
rect 67840 11450 67900 12420
rect 67840 10210 67900 11180
rect 67280 9940 67510 10130
rect 67990 11450 68050 12420
rect 67990 10210 68050 11180
rect 68150 11450 68210 12420
rect 68150 10210 68210 11180
rect 68310 11450 68370 12420
rect 68310 10210 68370 11180
rect 68860 12500 69090 12690
rect 68470 11450 68530 12420
rect 68470 10210 68530 11180
rect 67910 9940 68140 10130
rect 68630 11450 68690 12420
rect 68630 10210 68690 11180
rect 68780 11450 68840 12420
rect 68780 10210 68840 11180
rect 68940 11450 69000 12420
rect 68940 10210 69000 11180
rect 69490 12500 69720 12690
rect 69100 11450 69160 12420
rect 69100 10210 69160 11180
rect 68540 9940 68770 10130
rect 69260 11450 69320 12420
rect 69260 10210 69320 11180
rect 69420 11450 69480 12420
rect 69420 10210 69480 11180
rect 69580 11450 69640 12420
rect 69580 10210 69640 11180
rect 69730 11450 69790 12420
rect 69730 10210 69790 11180
rect 69180 9940 69400 10130
rect 69890 11450 69950 12420
rect 69890 10210 69950 11180
rect 70060 11450 70120 12420
rect 70060 10210 70120 11180
rect 69810 9940 70030 10130
rect 71210 9670 71580 9860
rect 71200 8710 71860 8910
rect 8220 7710 8900 8190
rect 12010 7710 12690 8190
rect 41190 7840 41560 8120
rect 42210 7840 42510 8120
rect 9110 6100 9250 7060
rect 9380 6100 9440 7060
rect 9540 6100 9600 7060
rect 9700 6100 9760 7060
rect 9890 6110 10030 7070
rect 12810 6100 12950 7060
rect 13080 6100 13140 7060
rect 13240 6100 13300 7060
rect 13400 6100 13460 7060
rect 13600 6100 13740 7060
rect 39240 6130 39410 7090
rect 8570 5130 8850 5310
rect 9110 4880 9250 5840
rect 9380 4880 9440 5840
rect 9540 4880 9600 5840
rect 9700 4880 9760 5840
rect 9890 4880 10030 5840
rect 12810 4880 12950 5840
rect 13080 4880 13140 5840
rect 13240 4880 13300 5840
rect 13400 4880 13460 5840
rect 13600 4880 13740 5840
rect 38630 5420 38860 6040
rect 39540 6130 39600 7090
rect 39690 6130 39750 7090
rect 39850 6130 39910 7090
rect 40010 6130 40070 7090
rect 40170 6130 40230 7090
rect 40330 6130 40390 7090
rect 40480 6130 40540 7090
rect 40640 6130 40700 7090
rect 40800 6130 40860 7090
rect 40960 6130 41020 7090
rect 41120 6130 41180 7090
rect 41270 6130 41330 7090
rect 41430 6130 41490 7090
rect 41590 6130 41650 7090
rect 41750 6130 41810 7090
rect 41940 6130 42110 7090
rect 44800 7030 45180 7410
rect 50730 7230 51280 7410
rect 46740 6410 47100 6790
rect 44200 5810 44580 6190
rect 47640 6130 47810 7090
rect 13970 5130 14250 5310
rect 47940 6130 48000 7090
rect 48090 6130 48150 7090
rect 48250 6130 48310 7090
rect 48410 6130 48470 7090
rect 48570 6130 48630 7090
rect 48730 6130 48790 7090
rect 48880 6130 48940 7090
rect 49040 6130 49100 7090
rect 49200 6130 49260 7090
rect 49360 6130 49420 7090
rect 49520 6130 49580 7090
rect 49670 6130 49730 7090
rect 49830 6130 49890 7090
rect 49990 6130 50050 7090
rect 50150 6130 50210 7090
rect 50340 6130 50510 7090
rect 81920 8350 82300 8590
rect 71200 8100 71860 8300
rect 66860 6940 66920 7900
rect 67120 6940 67180 7900
rect 67380 6940 67440 7900
rect 67640 6940 67700 7900
rect 67890 6940 67950 7900
rect 68150 6940 68210 7900
rect 68410 6940 68470 7900
rect 68670 6940 68730 7900
rect 68920 6940 68980 7900
rect 69180 6940 69240 7900
rect 69440 6940 69500 7900
rect 69700 6940 69760 7900
rect 69960 6940 70020 7900
rect 70220 6940 70280 7900
rect 70460 6940 70520 7900
rect 70720 6940 70780 7900
rect 70980 6940 71040 7900
rect 71240 6940 71300 7900
rect 71500 6940 71560 7900
rect 71760 6940 71820 7900
rect 72010 6940 72070 7900
rect 72270 6940 72330 7900
rect 72530 6940 72590 7900
rect 72790 6940 72850 7900
rect 73050 6940 73110 7900
rect 73310 6940 73370 7900
rect 73570 6940 73630 7900
rect 84250 6870 84310 7820
rect 84400 6870 84460 7820
rect 84560 6870 84620 7820
rect 84720 6870 84780 7820
rect 84880 6870 84940 7820
rect 85030 6870 85090 7820
rect 85190 6870 85250 7820
rect 85350 6870 85410 7820
rect 85510 6870 85570 7820
rect 85670 6870 85730 7820
rect 85820 6870 85880 7820
rect 85980 6870 86040 7820
rect 86140 6870 86200 7820
rect 50720 5810 51270 5990
rect 52530 5920 53290 6320
rect 66860 5700 66920 6660
rect 67120 5700 67180 6660
rect 67380 5700 67440 6660
rect 67640 5700 67700 6660
rect 67890 5700 67950 6660
rect 68150 5700 68210 6660
rect 68410 5700 68470 6660
rect 68670 5700 68730 6660
rect 68920 5700 68980 6660
rect 69180 5700 69240 6660
rect 69440 5700 69500 6660
rect 69700 5700 69760 6660
rect 69960 5700 70020 6660
rect 70220 5700 70280 6660
rect 70460 5700 70520 6660
rect 70720 5700 70780 6660
rect 70980 5700 71040 6660
rect 71240 5700 71300 6660
rect 71500 5700 71560 6660
rect 71760 5700 71820 6660
rect 72010 5700 72070 6660
rect 72270 5700 72330 6660
rect 72530 5700 72590 6660
rect 72790 5700 72850 6660
rect 73050 5700 73110 6660
rect 73310 5700 73370 6660
rect 83770 6670 84000 6780
rect 73570 5700 73630 6660
rect 84670 6670 84830 6780
rect 84250 5630 84310 6580
rect 84400 5630 84460 6580
rect 84560 5630 84620 6580
rect 84720 5630 84780 6580
rect 84880 5630 84940 6580
rect 85030 5630 85090 6580
rect 85190 5630 85250 6580
rect 85350 5630 85410 6580
rect 85510 5630 85570 6580
rect 85670 5630 85730 6580
rect 85820 5630 85880 6580
rect 85980 5630 86040 6580
rect 86140 5630 86200 6580
rect 47490 5100 47790 5280
rect 38770 3310 38830 3690
rect 39030 3310 39090 3690
rect 39290 3310 39350 4250
rect 39540 3310 39600 3690
rect 39800 3310 39860 4250
rect 40060 3310 40120 3690
rect 40320 3310 40380 4240
rect 40580 3310 40640 3690
rect 40830 3310 40890 4250
rect 41090 3310 41150 3690
rect 41350 3310 41410 4250
rect 41610 3310 41670 3690
rect 41870 3310 41930 4250
rect 42120 3310 42180 3690
rect 42380 3310 42440 4250
rect 42640 3310 42700 3690
rect 42900 3310 42960 4250
rect 43160 3310 43220 3690
rect 43410 3310 43470 4250
rect 43670 3310 43730 3690
rect 43930 3310 43990 4250
rect 44190 3310 44250 3690
rect 44450 3310 44510 4250
rect 44700 3310 44760 3690
rect 44960 3310 45020 4250
rect 45220 3310 45280 3690
rect 45480 3310 45540 4250
rect 45740 3310 45800 3690
rect 45990 3310 46050 3690
rect 39100 3110 39240 3230
rect 39400 3110 39750 3230
rect 39910 3110 40260 3230
rect 40430 3110 40780 3230
rect 40940 3110 41290 3230
rect 41460 3110 41810 3230
rect 41980 3110 42330 3230
rect 42490 3110 42840 3230
rect 43010 3110 43360 3230
rect 43520 3110 43870 3230
rect 44040 3110 44390 3230
rect 44560 3110 44910 3230
rect 45070 3110 45420 3230
rect 45590 3110 45730 3230
rect 38770 2090 38830 2470
rect 39030 2090 39090 2470
rect 39290 2090 39350 3030
rect 39540 2090 39600 2470
rect 39800 2090 39860 3030
rect 40060 2090 40120 2470
rect 40320 2090 40380 3030
rect 40580 2090 40640 2470
rect 40830 2090 40890 3030
rect 41090 2090 41150 2470
rect 41610 2090 41670 2470
rect 41870 2090 41930 3030
rect 42120 2090 42180 2470
rect 42380 2090 42440 3030
rect 42640 2090 42700 2470
rect 42900 2090 42960 3030
rect 43160 2090 43220 2470
rect 43410 2090 43470 3030
rect 43670 2090 43730 2470
rect 43930 2090 43990 3030
rect 44190 2090 44250 2470
rect 44450 2090 44510 3030
rect 44700 2090 44760 2470
rect 44960 2090 45020 3030
rect 45220 2090 45280 2470
rect 45480 2090 45540 3030
rect 47150 3250 47210 4210
rect 47420 3250 47480 4210
rect 45740 2090 45800 2470
rect 45990 2090 46050 2470
rect 47150 2020 47210 2980
rect 47670 3250 47730 4210
rect 47420 2020 47480 2980
rect 47670 2020 47730 2980
rect 47930 3250 47990 4210
rect 47930 2020 47990 2980
rect 48190 3250 48250 4210
rect 48450 3250 48510 4210
rect 48190 2020 48250 2980
rect 48700 3250 48760 4210
rect 48450 2020 48510 2980
rect 48700 2020 48760 2980
rect 48960 3250 49020 4210
rect 48960 2020 49020 2980
rect 49220 3250 49280 4210
rect 49480 3250 49540 4210
rect 49220 2020 49280 2980
rect 49740 3250 49800 4210
rect 49480 2020 49540 2980
rect 49740 2020 49800 2980
rect 49990 3250 50050 4210
rect 49990 2020 50050 2980
rect 50260 3250 50320 4210
rect 51010 4070 51230 4460
rect 66860 4460 66920 5420
rect 67120 4460 67180 5420
rect 67380 4460 67440 5420
rect 67640 4460 67700 5420
rect 67890 4460 67950 5420
rect 68150 4460 68210 5420
rect 68410 4460 68470 5420
rect 68670 4460 68730 5420
rect 68920 4460 68980 5420
rect 69180 4460 69240 5420
rect 69440 4460 69500 5420
rect 69700 4460 69760 5420
rect 69960 4460 70020 5420
rect 70220 4460 70280 5420
rect 70460 4460 70520 5420
rect 70720 4460 70780 5420
rect 70980 4460 71040 5420
rect 71240 4460 71300 5420
rect 71500 4460 71560 5420
rect 71760 4460 71820 5420
rect 72010 4460 72070 5420
rect 72270 4460 72330 5420
rect 72530 4460 72590 5420
rect 72790 4460 72850 5420
rect 73050 4460 73110 5420
rect 73310 4460 73370 5420
rect 73570 4460 73630 5420
rect 66860 3220 66920 4180
rect 67120 3220 67180 4180
rect 67380 3220 67440 4180
rect 67640 3220 67700 4180
rect 67890 3220 67950 4180
rect 68150 3220 68210 4180
rect 68410 3220 68470 4180
rect 68670 3220 68730 4180
rect 68920 3220 68980 4180
rect 69180 3220 69240 4180
rect 69440 3220 69500 4180
rect 69700 3220 69760 4180
rect 69960 3220 70020 4180
rect 70220 3220 70280 4180
rect 70460 3220 70520 4180
rect 70720 3220 70780 4180
rect 70980 3220 71040 4180
rect 71240 3220 71300 4180
rect 71500 3220 71560 4180
rect 71760 3220 71820 4180
rect 72010 3220 72070 4180
rect 72270 3220 72330 4180
rect 72530 3220 72590 4180
rect 72790 3220 72850 4180
rect 73050 3220 73110 4180
rect 73310 3220 73370 4180
rect 73570 3220 73630 4180
rect 84240 3540 84300 4490
rect 84390 3540 84450 4490
rect 84550 3540 84610 4490
rect 84710 3540 84770 4490
rect 84870 3540 84930 4490
rect 85020 3540 85080 4490
rect 85180 3540 85240 4490
rect 85340 3540 85400 4490
rect 85500 3540 85560 4490
rect 85660 3540 85720 4490
rect 85810 3540 85870 4490
rect 85970 3540 86030 4490
rect 86130 3540 86190 4490
rect 50260 2020 50320 2980
rect 84240 2310 84300 3260
rect 84390 2310 84450 3260
rect 84550 2310 84610 3260
rect 84710 2310 84770 3260
rect 84870 2310 84930 3260
rect 85020 2310 85080 3260
rect 85180 2310 85240 3260
rect 85340 2310 85400 3260
rect 85500 2310 85560 3260
rect 85660 2310 85720 3260
rect 85810 2310 85870 3260
rect 85970 2310 86030 3260
rect 86130 2310 86190 3260
rect 93240 2870 93620 3260
rect 51360 710 51590 920
rect 51790 850 52040 1010
rect 52190 900 52420 960
rect 53400 840 53620 1030
rect 7190 10 8770 390
<< metal2 >>
rect 2990 45140 3090 45150
rect 2990 44840 3000 45140
rect 3080 44840 3090 45140
rect 2990 44830 3090 44840
rect 3540 45140 3640 45150
rect 3540 44840 3550 45140
rect 3630 44840 3640 45140
rect 3540 44830 3640 44840
rect 4100 45140 4200 45150
rect 4100 44840 4110 45140
rect 4190 44840 4200 45140
rect 4100 44830 4200 44840
rect 4650 45140 4750 45150
rect 4650 44840 4660 45140
rect 4740 44840 4750 45140
rect 4650 44830 4750 44840
rect 5200 45140 5300 45150
rect 5200 44840 5210 45140
rect 5290 44840 5300 45140
rect 5200 44830 5300 44840
rect 5760 45140 5860 45150
rect 5760 44840 5770 45140
rect 5850 44840 5860 45140
rect 5760 44830 5860 44840
rect 6310 45140 6410 45150
rect 6310 44840 6320 45140
rect 6400 44840 6410 45140
rect 6310 44830 6410 44840
rect 6860 45140 6960 45150
rect 6860 44840 6870 45140
rect 6950 44840 6960 45140
rect 6860 44830 6960 44840
rect 7400 45140 7500 45150
rect 7400 44840 7410 45140
rect 7490 44840 7500 45140
rect 7400 44830 7500 44840
rect 7960 45140 8060 45150
rect 7960 44840 7970 45140
rect 8050 44840 8060 45140
rect 7960 44830 8060 44840
rect 8500 45140 8600 45150
rect 8500 44840 8510 45140
rect 8590 44840 8600 45140
rect 8500 44830 8600 44840
rect 9060 45140 9160 45150
rect 9060 44840 9070 45140
rect 9150 44840 9160 45140
rect 9060 44830 9160 44840
rect 9610 45140 9710 45150
rect 9610 44840 9620 45140
rect 9700 44840 9710 45140
rect 9610 44830 9710 44840
rect 10170 45140 10270 45150
rect 10170 44840 10180 45140
rect 10260 44840 10270 45140
rect 10170 44830 10270 44840
rect 10720 45140 10820 45150
rect 10720 44840 10730 45140
rect 10810 44840 10820 45140
rect 10720 44830 10820 44840
rect 11280 45140 11380 45150
rect 11280 44840 11290 45140
rect 11370 44840 11380 45140
rect 12380 45140 12480 45150
rect 11280 44830 11380 44840
rect 11880 44960 12150 44970
rect 11880 44770 11890 44960
rect 12140 44770 12150 44960
rect 12380 44840 12390 45140
rect 12470 44840 12480 45140
rect 12380 44830 12480 44840
rect 12930 45140 13030 45150
rect 12930 44840 12940 45140
rect 13020 44840 13030 45140
rect 12930 44830 13030 44840
rect 13470 45140 13570 45150
rect 13470 44840 13480 45140
rect 13560 44840 13570 45140
rect 13470 44830 13570 44840
rect 14030 45140 14130 45150
rect 14030 44840 14040 45140
rect 14120 44840 14130 45140
rect 14030 44830 14130 44840
rect 14580 45140 14680 45150
rect 14580 44840 14590 45140
rect 14670 44840 14680 45140
rect 14580 44830 14680 44840
rect 15130 45140 15230 45150
rect 15130 44840 15140 45140
rect 15220 44840 15230 45140
rect 15130 44830 15230 44840
rect 16240 45140 16340 45150
rect 16240 44840 16250 45140
rect 16330 44840 16340 45140
rect 16240 44830 16340 44840
rect 16790 45140 16890 45150
rect 16790 44840 16800 45140
rect 16880 44840 16890 45140
rect 16790 44830 16890 44840
rect 17340 45140 17440 45150
rect 17340 44840 17350 45140
rect 17430 44840 17440 45140
rect 17340 44830 17440 44840
rect 17900 45140 18000 45150
rect 17900 44840 17910 45140
rect 17990 44840 18000 45140
rect 17900 44830 18000 44840
rect 18450 45140 18550 45150
rect 18450 44840 18460 45140
rect 18540 44840 18550 45140
rect 18450 44830 18550 44840
rect 19000 45140 19100 45150
rect 19000 44840 19010 45140
rect 19090 44840 19100 45140
rect 19000 44830 19100 44840
rect 19550 45140 19650 45150
rect 19550 44840 19560 45140
rect 19640 44840 19650 45140
rect 19550 44830 19650 44840
rect 20110 45140 20210 45150
rect 20110 44840 20120 45140
rect 20200 44840 20210 45140
rect 20110 44830 20210 44840
rect 20660 45140 20760 45150
rect 20660 44840 20670 45140
rect 20750 44840 20760 45140
rect 20660 44830 20760 44840
rect 21210 45140 21310 45150
rect 21210 44840 21220 45140
rect 21300 44840 21310 45140
rect 21210 44830 21310 44840
rect 21760 45140 21860 45150
rect 21760 44840 21770 45140
rect 21850 44840 21860 45140
rect 21760 44830 21860 44840
rect 22300 45140 22400 45150
rect 22300 44840 22310 45140
rect 22390 44840 22400 45140
rect 22300 44830 22400 44840
rect 23360 45140 23550 45150
rect 23360 44960 23370 45140
rect 23540 44960 23550 45140
rect 11880 44760 12150 44770
rect 3500 44580 3650 44590
rect 3500 44440 3510 44580
rect 3640 44440 3650 44580
rect 3500 44430 3650 44440
rect 3510 43420 3640 44430
rect 23360 44040 23550 44960
rect 23970 45140 24070 45150
rect 23970 44840 23980 45140
rect 24060 44840 24070 45140
rect 24470 45140 24660 45150
rect 24470 44960 24480 45140
rect 24650 44960 24660 45140
rect 24470 44950 24660 44960
rect 25570 45140 25760 45150
rect 25570 44960 25580 45140
rect 25750 44960 25760 45140
rect 25570 44950 25760 44960
rect 27000 45010 27220 45020
rect 27000 44870 27010 45010
rect 27210 44870 27220 45010
rect 27000 44860 27220 44870
rect 23970 44830 24070 44840
rect 97760 44770 97940 44780
rect 97760 44630 97770 44770
rect 97930 44630 97940 44770
rect 23360 43960 23370 44040
rect 23540 43960 23550 44040
rect 23360 43950 23550 43960
rect 28100 44620 28370 44630
rect 97760 44620 97940 44630
rect 28100 44450 28110 44620
rect 28360 44450 28370 44620
rect 28100 43860 28370 44450
rect 28100 43700 28110 43860
rect 28360 43700 28370 43860
rect 28100 43690 28370 43700
rect 97850 43670 97940 44620
rect 97850 43580 98070 43670
rect 97980 43430 98070 43580
rect 70600 12960 70990 12970
rect 70600 12770 70610 12960
rect 70980 12770 70990 12960
rect 70600 12760 70990 12770
rect 66320 12690 66570 12700
rect 66320 12500 66330 12690
rect 66560 12500 66570 12690
rect 66320 12490 66570 12500
rect 66950 12690 67200 12700
rect 66950 12500 66960 12690
rect 67190 12500 67200 12690
rect 66950 12490 67200 12500
rect 67590 12690 67840 12700
rect 67590 12500 67600 12690
rect 67830 12500 67840 12690
rect 67590 12490 67840 12500
rect 68220 12690 68470 12700
rect 68220 12500 68230 12690
rect 68460 12500 68470 12690
rect 68220 12490 68470 12500
rect 68850 12690 69100 12700
rect 68850 12500 68860 12690
rect 69090 12500 69100 12690
rect 68850 12490 69100 12500
rect 69480 12690 69730 12700
rect 69480 12500 69490 12690
rect 69720 12500 69730 12690
rect 69480 12490 69730 12500
rect 66230 12420 66330 12430
rect 66230 11450 66250 12420
rect 66310 11450 66330 12420
rect 66230 11180 66330 11450
rect 66230 10790 66250 11180
rect 66310 10790 66330 11180
rect 66230 10410 66240 10790
rect 66320 10410 66330 10790
rect 66230 10210 66250 10410
rect 66310 10210 66330 10410
rect 66230 10200 66330 10210
rect 66400 12420 66490 12430
rect 66400 12080 66420 12420
rect 66400 11700 66410 12080
rect 66400 11450 66420 11700
rect 66480 11450 66490 12420
rect 66400 11180 66490 11450
rect 66400 10210 66420 11180
rect 66480 10210 66490 11180
rect 66400 10200 66490 10210
rect 66560 12420 66650 12430
rect 66560 11450 66570 12420
rect 66630 11450 66650 12420
rect 66560 11180 66650 11450
rect 66560 10210 66570 11180
rect 66630 10210 66650 11180
rect 66560 10200 66650 10210
rect 66720 12420 66810 12430
rect 66720 11450 66730 12420
rect 66790 11450 66810 12420
rect 66720 11430 66810 11450
rect 66720 10210 66730 11430
rect 66790 10210 66810 11430
rect 66720 10200 66810 10210
rect 66880 12420 66960 12430
rect 66880 11450 66890 12420
rect 66950 11450 66960 12420
rect 66880 11180 66960 11450
rect 66880 10210 66890 11180
rect 66950 10210 66960 11180
rect 66880 10200 66960 10210
rect 67030 12420 67120 12430
rect 67030 12080 67050 12420
rect 67030 11700 67040 12080
rect 67030 11450 67050 11700
rect 67110 11450 67120 12420
rect 67030 11180 67120 11450
rect 67030 10210 67050 11180
rect 67110 10210 67120 11180
rect 67030 10200 67120 10210
rect 67190 12420 67280 12430
rect 67190 11450 67200 12420
rect 67260 11450 67280 12420
rect 67190 11180 67280 11450
rect 67190 10210 67200 11180
rect 67260 10210 67280 11180
rect 67190 10200 67280 10210
rect 67350 12420 67440 12430
rect 67350 11450 67360 12420
rect 67420 11450 67440 12420
rect 67350 11430 67440 11450
rect 67350 10210 67360 11430
rect 67420 10210 67440 11430
rect 67350 10200 67440 10210
rect 67510 12420 67600 12430
rect 67510 11450 67520 12420
rect 67580 11450 67600 12420
rect 67510 11180 67600 11450
rect 67510 10210 67520 11180
rect 67580 10210 67600 11180
rect 67510 10200 67600 10210
rect 67670 12420 67750 12430
rect 67670 11450 67680 12420
rect 67740 11450 67750 12420
rect 67670 11180 67750 11450
rect 67670 10210 67680 11180
rect 67740 10210 67750 11180
rect 67670 10200 67750 10210
rect 67820 12420 67910 12430
rect 67820 11450 67840 12420
rect 67900 11450 67910 12420
rect 67820 11180 67910 11450
rect 67820 10210 67840 11180
rect 67900 10210 67910 11180
rect 67820 10200 67910 10210
rect 67980 12420 68070 12430
rect 67980 11450 67990 12420
rect 68050 11450 68070 12420
rect 67980 11430 68070 11450
rect 67980 10210 67990 11430
rect 68050 10210 68070 11430
rect 67980 10200 68070 10210
rect 68140 12420 68230 12430
rect 68140 11450 68150 12420
rect 68210 11450 68230 12420
rect 68140 11180 68230 11450
rect 68140 10210 68150 11180
rect 68210 10210 68230 11180
rect 68140 10200 68230 10210
rect 68300 12420 68390 12430
rect 68300 11450 68310 12420
rect 68370 12080 68390 12420
rect 68380 11700 68390 12080
rect 68370 11450 68390 11700
rect 68300 11180 68390 11450
rect 68300 10210 68310 11180
rect 68370 10210 68390 11180
rect 68300 10200 68390 10210
rect 68460 12420 68540 12430
rect 68460 11450 68470 12420
rect 68530 11450 68540 12420
rect 68460 11180 68540 11450
rect 68460 10210 68470 11180
rect 68530 10210 68540 11180
rect 68460 10200 68540 10210
rect 68610 12420 68700 12430
rect 68610 11450 68630 12420
rect 68690 11450 68700 12420
rect 68610 11430 68700 11450
rect 68610 11050 68620 11430
rect 68680 11180 68700 11430
rect 68610 10210 68630 11050
rect 68690 10210 68700 11180
rect 68610 10200 68700 10210
rect 68770 12420 68860 12430
rect 68770 11450 68780 12420
rect 68840 11450 68860 12420
rect 68770 11180 68860 11450
rect 68770 10210 68780 11180
rect 68840 10210 68860 11180
rect 68770 10200 68860 10210
rect 68930 12420 69020 12430
rect 68930 11450 68940 12420
rect 69000 12080 69020 12420
rect 69010 11700 69020 12080
rect 69000 11450 69020 11700
rect 68930 11180 69020 11450
rect 68930 10210 68940 11180
rect 69000 10210 69020 11180
rect 68930 10200 69020 10210
rect 69090 12420 69170 12430
rect 69090 11450 69100 12420
rect 69160 11450 69170 12420
rect 69090 11180 69170 11450
rect 69090 10210 69100 11180
rect 69160 10210 69170 11180
rect 69090 10200 69170 10210
rect 69240 12420 69330 12430
rect 69240 11450 69260 12420
rect 69320 11450 69330 12420
rect 69240 11430 69330 11450
rect 69240 11050 69250 11430
rect 69310 11180 69330 11430
rect 69240 10210 69260 11050
rect 69320 10210 69330 11180
rect 69240 10200 69330 10210
rect 69400 12420 69490 12430
rect 69400 11450 69420 12420
rect 69480 11450 69490 12420
rect 69400 11180 69490 11450
rect 69400 10210 69420 11180
rect 69480 10210 69490 11180
rect 69400 10200 69490 10210
rect 69560 12420 69650 12430
rect 69560 12080 69580 12420
rect 69560 11700 69570 12080
rect 69560 11450 69580 11700
rect 69640 11450 69650 12420
rect 69560 11180 69650 11450
rect 69560 10210 69580 11180
rect 69640 10210 69650 11180
rect 69560 10200 69650 10210
rect 69720 12420 69810 12430
rect 69720 11450 69730 12420
rect 69790 11450 69810 12420
rect 69720 11180 69810 11450
rect 69720 10210 69730 11180
rect 69790 10210 69810 11180
rect 69720 10200 69810 10210
rect 69880 12420 69970 12430
rect 69880 11450 69890 12420
rect 69950 11450 69970 12420
rect 69880 11430 69970 11450
rect 69880 10210 69890 11430
rect 69950 10210 69970 11430
rect 69880 10200 69970 10210
rect 70040 12420 70150 12430
rect 70040 11450 70060 12420
rect 70120 11450 70150 12420
rect 70040 11180 70150 11450
rect 70040 10210 70060 11180
rect 70120 10800 70150 11180
rect 70120 10400 71930 10800
rect 70120 10210 70150 10400
rect 70040 10200 70150 10210
rect 66640 10130 66880 10140
rect 53000 10090 53290 10100
rect 15740 9330 16400 9340
rect 3380 9250 3860 9260
rect 3380 8710 3390 9250
rect 3850 8710 3860 9250
rect 15740 8970 15750 9330
rect 16390 8970 16400 9330
rect 15740 8960 16400 8970
rect 19510 9320 19990 9330
rect 12950 8900 13220 8910
rect 3380 8700 3860 8710
rect 9250 8890 9520 8900
rect 9250 8580 9260 8890
rect 9510 8580 9520 8890
rect 9250 8570 9520 8580
rect 9620 8890 9890 8900
rect 9620 8580 9630 8890
rect 9880 8580 9890 8890
rect 12950 8590 12960 8900
rect 13210 8590 13220 8900
rect 12950 8580 13220 8590
rect 13320 8900 13590 8910
rect 13320 8590 13330 8900
rect 13580 8590 13590 8900
rect 19510 8780 19520 9320
rect 19980 8780 19990 9320
rect 19510 8770 19990 8780
rect 27650 8790 30240 8860
rect 27650 8780 30310 8790
rect 13320 8580 13590 8590
rect 27650 8610 29720 8780
rect 9620 8570 9890 8580
rect 8200 8190 8920 8200
rect 8200 7710 8220 8190
rect 8900 7710 8920 8190
rect 8200 7700 8920 7710
rect 9100 7060 9260 7070
rect 9100 6100 9110 7060
rect 9250 6100 9260 7060
rect 9100 6090 9260 6100
rect 9370 7060 9450 8570
rect 9370 6100 9380 7060
rect 9440 6100 9450 7060
rect 9370 6090 9450 6100
rect 9530 7060 9610 7070
rect 9530 6100 9540 7060
rect 9600 6100 9610 7060
rect 9530 6090 9610 6100
rect 9690 7060 9770 8570
rect 12000 8190 12700 8200
rect 12000 7710 12010 8190
rect 12690 7710 12700 8190
rect 12000 7700 12700 7710
rect 9690 6100 9700 7060
rect 9760 6100 9770 7060
rect 9880 7070 10040 7080
rect 9880 6110 9890 7070
rect 10030 6110 10040 7070
rect 9880 6100 10040 6110
rect 12800 7060 12960 7070
rect 12800 6100 12810 7060
rect 12950 6100 12960 7060
rect 9100 5840 9260 5850
rect 8560 5310 8860 5320
rect 8560 5130 8570 5310
rect 8850 5130 8860 5310
rect 8560 5120 8860 5130
rect 9100 4880 9110 5840
rect 9250 4880 9260 5840
rect 9100 4870 9260 4880
rect 9370 5840 9450 5850
rect 9370 4880 9380 5840
rect 9440 4880 9450 5840
rect 9370 4870 9450 4880
rect 9530 5840 9610 5850
rect 9530 4880 9540 5840
rect 9600 4880 9610 5840
rect 9530 4870 9610 4880
rect 9690 5840 9770 6100
rect 12800 6090 12960 6100
rect 13070 7060 13150 8580
rect 13070 6100 13080 7060
rect 13140 6100 13150 7060
rect 9690 4880 9700 5840
rect 9760 4880 9770 5840
rect 9690 4870 9770 4880
rect 9880 5840 10040 5850
rect 9880 4880 9890 5840
rect 10030 4880 10040 5840
rect 9880 4870 10040 4880
rect 12800 5840 12960 5850
rect 12800 4880 12810 5840
rect 12950 4880 12960 5840
rect 12800 4870 12960 4880
rect 13070 5840 13150 6100
rect 13230 7060 13310 7070
rect 13230 6100 13240 7060
rect 13300 6100 13310 7060
rect 13230 6090 13310 6100
rect 13390 7060 13470 8580
rect 27650 8390 28700 8610
rect 27650 7430 27940 8390
rect 29080 8190 29720 8610
rect 30300 8190 30310 8780
rect 29080 8180 30310 8190
rect 13390 6100 13400 7060
rect 13460 6100 13470 7060
rect 13390 6090 13470 6100
rect 13590 7060 13750 7070
rect 13590 6100 13600 7060
rect 13740 6100 13750 7060
rect 27650 7030 28630 7430
rect 37970 6800 38250 9620
rect 41180 8120 41570 9560
rect 41180 7840 41190 8120
rect 41560 7840 41570 8120
rect 41180 7830 41570 7840
rect 41740 7700 42030 9880
rect 53000 9490 53010 10090
rect 53280 9490 53290 10090
rect 66640 9940 66650 10130
rect 66870 9940 66880 10130
rect 66640 9930 66880 9940
rect 67270 10130 67520 10140
rect 67270 9940 67280 10130
rect 67510 9940 67520 10130
rect 67270 9930 67520 9940
rect 67900 10130 68150 10140
rect 67900 9940 67910 10130
rect 68140 9940 68150 10130
rect 67900 9930 68150 9940
rect 68530 10130 68780 10140
rect 68530 9940 68540 10130
rect 68770 9940 68780 10130
rect 68530 9930 68780 9940
rect 69170 10130 69410 10140
rect 69170 9940 69180 10130
rect 69400 9940 69410 10130
rect 69170 9930 69410 9940
rect 69800 10130 70040 10140
rect 69800 9940 69810 10130
rect 70030 9940 70040 10130
rect 69800 9930 70040 9940
rect 53000 9480 53290 9490
rect 42200 8120 42520 8130
rect 42200 7840 42210 8120
rect 42510 7840 42520 8120
rect 42200 7830 42520 7840
rect 41740 7520 42130 7700
rect 39440 7450 41660 7460
rect 39440 7270 39450 7450
rect 41650 7270 41660 7450
rect 39440 7260 41660 7270
rect 39230 7090 39420 7100
rect 37950 6790 38280 6800
rect 37950 6410 37960 6790
rect 38270 6410 38280 6790
rect 37950 6400 38280 6410
rect 39230 6130 39240 7090
rect 39410 6130 39420 7090
rect 39230 6120 39420 6130
rect 39530 7090 39610 7260
rect 39530 6130 39540 7090
rect 39600 6130 39610 7090
rect 39530 6120 39610 6130
rect 39680 7090 39760 7100
rect 39680 6130 39690 7090
rect 39750 6130 39760 7090
rect 39680 6120 39760 6130
rect 39840 7090 39920 7100
rect 39840 6130 39850 7090
rect 39910 6130 39920 7090
rect 13590 6090 13750 6100
rect 38620 6040 38870 6050
rect 13070 4880 13080 5840
rect 13140 4880 13150 5840
rect 13070 4870 13150 4880
rect 13230 5840 13310 5850
rect 13230 4880 13240 5840
rect 13300 4880 13310 5840
rect 13230 4870 13310 4880
rect 13390 5840 13470 5850
rect 13390 4810 13400 5840
rect 13460 4810 13470 5840
rect 13590 5840 13750 5850
rect 13590 4880 13600 5840
rect 13740 4880 13750 5840
rect 38620 5420 38630 6040
rect 38860 5420 38870 6040
rect 39840 5950 39920 6130
rect 40000 7090 40080 7100
rect 40000 6130 40010 7090
rect 40070 6130 40080 7090
rect 40000 6120 40080 6130
rect 40160 7090 40240 7260
rect 40160 6130 40170 7090
rect 40230 6130 40240 7090
rect 40160 6120 40240 6130
rect 40320 7090 40400 7100
rect 40320 6130 40330 7090
rect 40390 6130 40400 7090
rect 40320 6120 40400 6130
rect 40470 7090 40550 7100
rect 40470 6130 40480 7090
rect 40540 6130 40550 7090
rect 40470 5950 40550 6130
rect 40630 7090 40710 7100
rect 40630 6130 40640 7090
rect 40700 6130 40710 7090
rect 40630 6120 40710 6130
rect 40790 7090 40870 7260
rect 40790 6130 40800 7090
rect 40860 6130 40870 7090
rect 40790 6120 40870 6130
rect 40950 7090 41030 7100
rect 40950 6130 40960 7090
rect 41020 6130 41030 7090
rect 40950 6120 41030 6130
rect 41110 7090 41190 7100
rect 41110 6130 41120 7090
rect 41180 6130 41190 7090
rect 41110 5950 41190 6130
rect 41260 7090 41340 7100
rect 41260 6130 41270 7090
rect 41330 6130 41340 7090
rect 41260 6120 41340 6130
rect 41420 7090 41500 7260
rect 41420 6130 41430 7090
rect 41490 6130 41500 7090
rect 41420 6120 41500 6130
rect 41580 7090 41660 7100
rect 41580 6130 41590 7090
rect 41650 6130 41660 7090
rect 41580 6120 41660 6130
rect 41740 7090 41820 7100
rect 41740 6130 41750 7090
rect 41810 6130 41820 7090
rect 41740 5950 41820 6130
rect 39440 5940 41820 5950
rect 39440 5760 39450 5940
rect 41810 5760 41820 5940
rect 39440 5750 41820 5760
rect 41930 7090 42130 7520
rect 41930 6130 41940 7090
rect 42110 6130 42130 7090
rect 38620 5410 38870 5420
rect 13960 5310 14260 5320
rect 13960 5130 13970 5310
rect 14250 5130 14260 5310
rect 40760 5250 40960 5260
rect 13960 5120 14260 5130
rect 13590 4870 13750 4880
rect 13390 4800 13470 4810
rect 3000 1710 3840 4730
rect 6780 2860 7620 4720
rect 6780 2000 16240 2860
rect 3000 1700 12180 1710
rect 3000 830 12340 1700
rect 11340 490 12340 830
rect 7180 390 8780 400
rect 7180 10 7190 390
rect 8770 10 8780 390
rect 7180 0 8780 10
rect 11340 10 11350 490
rect 12330 10 12340 490
rect 11340 0 12340 10
rect 15240 490 16240 2000
rect 15240 10 15250 490
rect 16230 10 16240 490
rect 15240 0 16240 10
rect 18100 840 18960 4710
rect 21840 880 22700 4710
rect 25620 880 26480 4730
rect 27650 2660 28360 4720
rect 27640 2560 28360 2660
rect 27640 2550 28520 2560
rect 27640 2540 28660 2550
rect 27640 2320 27670 2540
rect 27660 2060 27670 2320
rect 28650 2060 28660 2540
rect 27660 2050 28660 2060
rect 33640 1960 34020 5200
rect 40760 4870 40770 5250
rect 40950 4870 40960 5250
rect 41930 4900 42130 6130
rect 40760 4860 40960 4870
rect 37410 4260 37800 4840
rect 39730 4720 39930 4730
rect 39730 4340 39740 4720
rect 39920 4340 39930 4720
rect 39730 4330 39930 4340
rect 37410 4250 39360 4260
rect 37410 3840 39290 4250
rect 38770 3690 38830 3700
rect 38770 3300 38830 3310
rect 39030 3690 39090 3700
rect 39030 3300 39090 3310
rect 39280 3310 39290 3840
rect 39350 3310 39360 4250
rect 39790 4250 39870 4330
rect 39280 3300 39360 3310
rect 39540 3690 39600 3700
rect 39540 3300 39600 3310
rect 39790 3310 39800 4250
rect 39860 3310 39870 4250
rect 40820 4250 40900 4860
rect 40250 4230 40320 4240
rect 40380 4230 40450 4240
rect 40250 3850 40260 4230
rect 40440 3850 40450 4230
rect 40250 3840 40320 3850
rect 39790 3300 39870 3310
rect 40060 3690 40120 3700
rect 40060 3300 40120 3310
rect 40310 3310 40320 3840
rect 40380 3840 40450 3850
rect 40380 3310 40390 3840
rect 39090 3230 39250 3240
rect 39090 3110 39100 3230
rect 39240 3110 39250 3230
rect 39090 3100 39250 3110
rect 39390 3230 39760 3240
rect 39390 3110 39400 3230
rect 39750 3110 39760 3230
rect 39390 3100 39760 3110
rect 39900 3230 40270 3240
rect 39900 3110 39910 3230
rect 40260 3110 40270 3230
rect 39900 3100 40270 3110
rect 39280 3030 39360 3040
rect 39280 3000 39290 3030
rect 39220 2990 39290 3000
rect 39350 3000 39360 3030
rect 39790 3030 39870 3040
rect 39350 2990 39420 3000
rect 39220 2610 39230 2990
rect 39410 2610 39420 2990
rect 39220 2600 39290 2610
rect 38770 2470 38830 2480
rect 38770 2080 38830 2090
rect 39030 2470 39090 2480
rect 39030 2080 39090 2090
rect 39280 2090 39290 2600
rect 39350 2600 39420 2610
rect 39350 2090 39360 2600
rect 39280 2080 39360 2090
rect 39540 2470 39600 2480
rect 39540 2080 39600 2090
rect 39790 2090 39800 3030
rect 39860 2090 39870 3030
rect 40310 3030 40390 3310
rect 40580 3690 40640 3700
rect 40580 3300 40640 3310
rect 40820 3310 40830 4250
rect 40890 3310 40900 4250
rect 41340 4690 42130 4900
rect 41340 4250 41420 4690
rect 40420 3230 40790 3240
rect 40420 3110 40430 3230
rect 40780 3110 40790 3230
rect 40420 3100 40790 3110
rect 39790 1970 39870 2090
rect 40060 2470 40120 2480
rect 40060 2080 40120 2090
rect 40310 2090 40320 3030
rect 40380 2090 40390 3030
rect 40820 3030 40900 3310
rect 41090 3690 41150 3700
rect 41090 3300 41150 3310
rect 41340 3310 41350 4250
rect 41410 3310 41420 4250
rect 41860 4250 41940 4690
rect 42320 4260 42520 7830
rect 42830 4740 43030 9030
rect 44790 7410 45190 7420
rect 44790 7030 44800 7410
rect 45180 7030 45190 7410
rect 44790 7020 45190 7030
rect 45530 6790 45930 9350
rect 53450 8760 53840 9340
rect 51920 8470 53840 8760
rect 60100 8860 60440 9200
rect 64080 9080 69920 9460
rect 64400 8860 68360 8980
rect 60100 8600 68360 8860
rect 50720 7410 51290 7420
rect 50720 7230 50730 7410
rect 51280 7230 51290 7410
rect 50720 7220 51290 7230
rect 47630 7090 47820 7100
rect 45530 6410 45540 6790
rect 45920 6410 45930 6790
rect 45530 6400 45930 6410
rect 46730 6790 47110 6800
rect 46730 6410 46740 6790
rect 47100 6410 47110 6790
rect 46730 6400 47110 6410
rect 44190 6190 44590 6200
rect 44190 5810 44200 6190
rect 44580 5810 44590 6190
rect 47630 6130 47640 7090
rect 47810 6130 47820 7090
rect 47630 6120 47820 6130
rect 47930 7090 48010 7100
rect 47930 6130 47940 7090
rect 48000 6130 48010 7090
rect 47930 6080 48010 6130
rect 48080 7090 48160 7100
rect 48080 6130 48090 7090
rect 48150 6130 48160 7090
rect 48080 6120 48160 6130
rect 48240 7090 48320 7100
rect 48240 6130 48250 7090
rect 48310 6130 48320 7090
rect 48240 6080 48320 6130
rect 48400 7090 48480 7100
rect 48400 6130 48410 7090
rect 48470 6130 48480 7090
rect 48400 6120 48480 6130
rect 48560 7090 48640 7100
rect 48560 6130 48570 7090
rect 48630 6130 48640 7090
rect 48560 6080 48640 6130
rect 48720 7090 48800 7100
rect 48720 6130 48730 7090
rect 48790 6130 48800 7090
rect 48720 6120 48800 6130
rect 48870 7090 48950 7100
rect 48870 6130 48880 7090
rect 48940 6130 48950 7090
rect 48870 6080 48950 6130
rect 49030 7090 49110 7100
rect 49030 6130 49040 7090
rect 49100 6130 49110 7090
rect 49030 6120 49110 6130
rect 49190 7090 49270 7100
rect 49190 6130 49200 7090
rect 49260 6130 49270 7090
rect 49190 6080 49270 6130
rect 49350 7090 49430 7100
rect 49350 6130 49360 7090
rect 49420 6130 49430 7090
rect 49350 6120 49430 6130
rect 49510 7090 49590 7100
rect 49510 6130 49520 7090
rect 49580 6130 49590 7090
rect 49510 6080 49590 6130
rect 49660 7090 49740 7100
rect 49660 6130 49670 7090
rect 49730 6130 49740 7090
rect 49660 6120 49740 6130
rect 49820 7090 49900 7100
rect 49820 6130 49830 7090
rect 49890 6130 49900 7090
rect 49820 6080 49900 6130
rect 49980 7090 50060 7100
rect 49980 6130 49990 7090
rect 50050 6130 50060 7090
rect 49980 6120 50060 6130
rect 50140 7090 50220 7100
rect 50140 6130 50150 7090
rect 50210 6130 50220 7090
rect 50140 6080 50220 6130
rect 50330 7090 50530 7100
rect 50330 6130 50340 7090
rect 50510 6130 50530 7090
rect 50330 6120 50530 6130
rect 44190 5800 44590 5810
rect 47890 5680 48050 6080
rect 47890 5390 47900 5680
rect 48040 5390 48050 5680
rect 47890 5380 48050 5390
rect 43860 5280 44590 5290
rect 43860 5100 43870 5280
rect 44580 5100 44590 5280
rect 43860 5090 44590 5100
rect 47480 5280 47800 5290
rect 47480 5100 47490 5280
rect 47790 5100 47800 5280
rect 47480 5090 47800 5100
rect 48200 5140 48350 6080
rect 48520 5680 48680 6080
rect 48520 5390 48530 5680
rect 48670 5390 48680 5680
rect 48520 5380 48680 5390
rect 48830 5140 48980 6080
rect 49150 5680 49310 6080
rect 49150 5390 49160 5680
rect 49300 5390 49310 5680
rect 49150 5380 49310 5390
rect 49480 5140 49630 6080
rect 49780 5680 49940 6080
rect 49780 5390 49790 5680
rect 49930 5390 49940 5680
rect 49780 5380 49940 5390
rect 50100 5140 50250 6080
rect 50710 5990 51280 6000
rect 50710 5810 50720 5990
rect 51270 5810 51280 5990
rect 50710 5800 51280 5810
rect 42830 4540 43550 4740
rect 42830 4260 43030 4540
rect 41340 3300 41420 3310
rect 41610 3690 41670 3700
rect 41610 3300 41670 3310
rect 41860 3310 41870 4250
rect 41930 3310 41940 4250
rect 42370 4250 42450 4260
rect 41860 3300 41940 3310
rect 42120 3690 42180 3700
rect 42120 3300 42180 3310
rect 42370 3310 42380 4250
rect 42440 3310 42450 4250
rect 42890 4250 42970 4260
rect 43350 4250 43550 4540
rect 43860 4260 44060 5090
rect 44380 5010 45110 5020
rect 44380 4830 44390 5010
rect 45100 4830 45110 5010
rect 48200 4940 50250 5140
rect 51920 5230 52310 8470
rect 66280 7980 67750 8180
rect 68000 7980 68360 8600
rect 68620 8460 69280 8480
rect 68620 8080 68640 8460
rect 69260 8130 69280 8460
rect 69260 8080 69290 8130
rect 68620 7980 69290 8080
rect 69540 7980 69920 9080
rect 70280 8620 70500 10400
rect 71200 9860 71590 9870
rect 71200 9670 71210 9860
rect 71580 9670 71590 9860
rect 71200 9660 71590 9670
rect 71870 8920 72360 9350
rect 82950 8940 83420 9340
rect 71190 8910 72360 8920
rect 71190 8710 71200 8910
rect 71860 8710 72360 8910
rect 71190 8700 72360 8710
rect 70280 8360 75300 8620
rect 52520 6320 53300 6330
rect 66280 6320 66660 7980
rect 52520 5920 52530 6320
rect 53290 5920 53300 6320
rect 63820 5940 66660 6320
rect 66810 7900 66970 7910
rect 66810 6940 66860 7900
rect 66920 6940 66970 7900
rect 66810 6660 66970 6940
rect 67070 7900 67230 7980
rect 67070 6940 67120 7900
rect 67180 6940 67230 7900
rect 67070 6930 67230 6940
rect 67330 7900 67490 7910
rect 67330 6940 67380 7900
rect 67440 6940 67490 7900
rect 52520 5910 53300 5920
rect 44380 4820 45110 4830
rect 44380 4260 44580 4820
rect 44890 4740 45620 4750
rect 44890 4560 44900 4740
rect 45610 4560 45620 4740
rect 44890 4550 45620 4560
rect 44890 4260 45090 4550
rect 45410 4260 45610 4550
rect 43920 4250 44000 4260
rect 40930 3230 41300 3240
rect 40930 3110 40940 3230
rect 41290 3110 41300 3230
rect 40930 3100 41300 3110
rect 41450 3230 41820 3240
rect 41450 3110 41460 3230
rect 41810 3110 41820 3230
rect 41450 3100 41820 3110
rect 41970 3230 42340 3240
rect 41970 3110 41980 3230
rect 42330 3110 42340 3230
rect 41970 3100 42340 3110
rect 40310 2080 40390 2090
rect 40580 2470 40640 2480
rect 40580 2080 40640 2090
rect 40820 2090 40830 3030
rect 40890 2090 40900 3030
rect 41810 3030 41990 3040
rect 40820 2080 40900 2090
rect 41090 2470 41150 2480
rect 41090 2080 41150 2090
rect 41610 2470 41670 2480
rect 41610 2080 41670 2090
rect 41810 2090 41870 3030
rect 41930 2090 41990 3030
rect 42370 3030 42450 3310
rect 42640 3690 42700 3700
rect 42640 3300 42700 3310
rect 42890 3310 42900 4250
rect 42960 3310 42970 4250
rect 42480 3230 42850 3240
rect 42480 3110 42490 3230
rect 42840 3110 42850 3230
rect 42480 3100 42850 3110
rect 33640 1580 33650 1960
rect 34010 1580 34020 1960
rect 33640 1570 34020 1580
rect 39730 1960 39930 1970
rect 39730 1580 39740 1960
rect 39920 1580 39930 1960
rect 39730 1570 39930 1580
rect 41810 1640 41990 2090
rect 42120 2470 42180 2480
rect 42120 2080 42180 2090
rect 42370 2090 42380 3030
rect 42440 2090 42450 3030
rect 42890 3030 42970 3310
rect 43160 3690 43220 3700
rect 43160 3300 43220 3310
rect 43400 3310 43410 4250
rect 43470 3310 43480 4250
rect 43000 3230 43370 3240
rect 43000 3110 43010 3230
rect 43360 3110 43370 3230
rect 43000 3100 43370 3110
rect 42370 2080 42450 2090
rect 42640 2470 42700 2480
rect 42640 2080 42700 2090
rect 42890 2090 42900 3030
rect 42960 2090 42970 3030
rect 43400 3030 43480 3310
rect 43670 3690 43730 3700
rect 43670 3300 43730 3310
rect 43920 3310 43930 4250
rect 43990 3310 44000 4250
rect 44440 4250 44520 4260
rect 43510 3230 43880 3240
rect 43510 3110 43520 3230
rect 43870 3110 43880 3230
rect 43510 3100 43880 3110
rect 42890 2080 42970 2090
rect 43160 2470 43220 2480
rect 43160 2080 43220 2090
rect 43400 2090 43410 3030
rect 43470 2090 43480 3030
rect 43920 3030 44000 3310
rect 44190 3690 44250 3700
rect 44190 3300 44250 3310
rect 44440 3310 44450 4250
rect 44510 3310 44520 4250
rect 44950 4250 45030 4260
rect 44030 3230 44400 3240
rect 44030 3110 44040 3230
rect 44390 3110 44400 3230
rect 44030 3100 44400 3110
rect 43400 2080 43480 2090
rect 43670 2470 43730 2480
rect 43670 2080 43730 2090
rect 43920 2090 43930 3030
rect 43990 2090 44000 3030
rect 44440 3030 44520 3310
rect 44700 3690 44760 3700
rect 44700 3300 44760 3310
rect 44950 3310 44960 4250
rect 45020 3310 45030 4250
rect 45470 4250 45550 4260
rect 44550 3230 44920 3240
rect 44550 3110 44560 3230
rect 44910 3110 44920 3230
rect 44550 3100 44920 3110
rect 43920 2080 44000 2090
rect 44190 2470 44250 2480
rect 44190 2080 44250 2090
rect 44440 2090 44450 3030
rect 44510 2090 44520 3030
rect 44950 3030 45030 3310
rect 45220 3690 45280 3700
rect 45220 3300 45280 3310
rect 45470 3310 45480 4250
rect 45540 3310 45550 4250
rect 48390 4240 48570 4940
rect 49430 4250 49610 4940
rect 51920 4830 51930 5230
rect 52300 4830 52310 5230
rect 51920 4820 52310 4830
rect 66810 5700 66860 6660
rect 66920 5700 66970 6660
rect 66810 5420 66970 5700
rect 51000 4460 51240 4470
rect 47140 4210 47220 4220
rect 45060 3230 45430 3240
rect 45060 3110 45070 3230
rect 45420 3110 45430 3230
rect 45060 3100 45430 3110
rect 44440 2080 44520 2090
rect 44700 2470 44760 2480
rect 44700 2080 44760 2090
rect 44950 2090 44960 3030
rect 45020 2090 45030 3030
rect 45470 3030 45550 3310
rect 45740 3690 45800 3700
rect 45740 3300 45800 3310
rect 45990 3690 46050 3700
rect 47140 3640 47150 4210
rect 45990 3300 46050 3310
rect 47100 3630 47150 3640
rect 47210 3640 47220 4210
rect 47410 4210 47490 4220
rect 47210 3630 47260 3640
rect 47100 3250 47110 3630
rect 47250 3250 47260 3630
rect 47100 3240 47260 3250
rect 47410 3250 47420 4210
rect 47480 3250 47490 4210
rect 47660 4210 47740 4220
rect 47660 3640 47670 4210
rect 45580 3230 45740 3240
rect 45580 3110 45590 3230
rect 45730 3110 45740 3230
rect 45580 3100 45740 3110
rect 44950 2080 45030 2090
rect 45220 2470 45280 2480
rect 45220 2080 45280 2090
rect 45470 2090 45480 3030
rect 45540 2090 45550 3030
rect 47140 2980 47220 3240
rect 47410 3060 47490 3250
rect 47620 3630 47670 3640
rect 47730 3640 47740 4210
rect 47880 4210 48040 4220
rect 47880 3830 47890 4210
rect 48030 3830 48040 4210
rect 47880 3820 47930 3830
rect 47730 3630 47780 3640
rect 47620 3250 47630 3630
rect 47770 3250 47780 3630
rect 47620 3240 47780 3250
rect 47920 3250 47930 3820
rect 47990 3820 48040 3830
rect 48180 4210 48260 4220
rect 47990 3250 48000 3820
rect 48180 3640 48190 4210
rect 45470 2080 45550 2090
rect 45740 2470 45800 2480
rect 45740 2080 45800 2090
rect 45990 2470 46050 2480
rect 45990 2080 46050 2090
rect 47140 2020 47150 2980
rect 47210 2020 47220 2980
rect 47370 3050 47530 3060
rect 47370 2670 47380 3050
rect 47520 2670 47530 3050
rect 47370 2660 47420 2670
rect 47140 2010 47220 2020
rect 47410 2020 47420 2660
rect 47480 2660 47530 2670
rect 47660 2980 47740 3240
rect 47480 2020 47490 2660
rect 47410 2010 47490 2020
rect 47660 2020 47670 2980
rect 47730 2020 47740 2980
rect 47660 2010 47740 2020
rect 47920 2980 48000 3250
rect 48140 3630 48190 3640
rect 48250 3640 48260 4210
rect 48440 4210 48520 4240
rect 48250 3630 48300 3640
rect 48140 3250 48150 3630
rect 48290 3250 48300 3630
rect 48140 3240 48300 3250
rect 48440 3250 48450 4210
rect 48510 3250 48520 4210
rect 48690 4210 48770 4220
rect 48690 3640 48700 4210
rect 47920 2020 47930 2980
rect 47990 2020 48000 2980
rect 47920 2010 48000 2020
rect 48180 2980 48260 3240
rect 48440 3060 48520 3250
rect 48650 3630 48700 3640
rect 48760 3640 48770 4210
rect 48910 4210 49070 4220
rect 48910 3830 48920 4210
rect 49060 3830 49070 4210
rect 48910 3820 48960 3830
rect 48760 3630 48810 3640
rect 48650 3250 48660 3630
rect 48800 3250 48810 3630
rect 48650 3240 48810 3250
rect 48950 3250 48960 3820
rect 49020 3820 49070 3830
rect 49210 4210 49290 4220
rect 49020 3250 49030 3820
rect 49210 3640 49220 4210
rect 48180 2020 48190 2980
rect 48250 2020 48260 2980
rect 48400 3050 48560 3060
rect 48400 2670 48410 3050
rect 48550 2670 48560 3050
rect 48400 2660 48450 2670
rect 48180 2010 48260 2020
rect 48440 2020 48450 2660
rect 48510 2660 48560 2670
rect 48690 2980 48770 3240
rect 48510 2020 48520 2660
rect 48440 2010 48520 2020
rect 48690 2020 48700 2980
rect 48760 2020 48770 2980
rect 48690 2010 48770 2020
rect 48950 2980 49030 3250
rect 49170 3630 49220 3640
rect 49280 3640 49290 4210
rect 49470 4210 49550 4250
rect 49280 3630 49330 3640
rect 49170 3250 49180 3630
rect 49320 3250 49330 3630
rect 49170 3240 49330 3250
rect 49470 3250 49480 4210
rect 49540 3250 49550 4210
rect 49730 4210 49810 4220
rect 49730 3640 49740 4210
rect 48950 2020 48960 2980
rect 49020 2020 49030 2980
rect 48950 2010 49030 2020
rect 49210 2980 49290 3240
rect 49470 3060 49550 3250
rect 49690 3630 49740 3640
rect 49800 3640 49810 4210
rect 49940 4210 50100 4220
rect 49940 3830 49950 4210
rect 50090 3830 50100 4210
rect 49940 3820 49990 3830
rect 49800 3630 49850 3640
rect 49690 3250 49700 3630
rect 49840 3250 49850 3630
rect 49690 3240 49850 3250
rect 49980 3250 49990 3820
rect 50050 3820 50100 3830
rect 50250 4210 50330 4220
rect 50050 3250 50060 3820
rect 50250 3640 50260 4210
rect 49210 2020 49220 2980
rect 49280 2020 49290 2980
rect 49430 3050 49590 3060
rect 49430 2670 49440 3050
rect 49580 2670 49590 3050
rect 49430 2660 49480 2670
rect 49210 2010 49290 2020
rect 49470 2020 49480 2660
rect 49540 2660 49590 2670
rect 49730 2980 49810 3240
rect 49540 2020 49550 2660
rect 49470 2010 49550 2020
rect 49730 2020 49740 2980
rect 49800 2020 49810 2980
rect 49730 2010 49810 2020
rect 49980 2980 50060 3250
rect 50210 3630 50260 3640
rect 50320 3640 50330 4210
rect 51000 4070 51010 4460
rect 51230 4070 51240 4460
rect 51000 4060 51240 4070
rect 50320 3630 50370 3640
rect 50210 3250 50220 3630
rect 50360 3250 50370 3630
rect 50210 3240 50370 3250
rect 59280 3500 59680 3520
rect 49980 2020 49990 2980
rect 50050 2020 50060 2980
rect 49980 2010 50060 2020
rect 50250 2980 50330 3240
rect 50250 2020 50260 2980
rect 50320 2020 50330 2980
rect 59280 2860 59300 3500
rect 59660 2860 59680 3500
rect 59280 2660 59680 2860
rect 60040 3140 60440 4720
rect 66810 4460 66860 5420
rect 66920 4460 66970 5420
rect 66810 4180 66970 4460
rect 66810 3800 66860 4180
rect 66920 3800 66970 4180
rect 66810 3220 66820 3800
rect 66960 3220 66970 3800
rect 66810 3210 66970 3220
rect 67070 6660 67230 6670
rect 67070 5700 67120 6660
rect 67180 5700 67230 6660
rect 67070 5420 67230 5700
rect 67070 4460 67120 5420
rect 67180 4460 67230 5420
rect 67070 4180 67230 4460
rect 67070 3220 67120 4180
rect 67180 3220 67230 4180
rect 67070 3140 67230 3220
rect 67330 6660 67490 6940
rect 67330 5700 67380 6660
rect 67440 5700 67490 6660
rect 67330 5420 67490 5700
rect 67590 7900 67750 7980
rect 67590 6940 67640 7900
rect 67700 6940 67750 7900
rect 67590 6660 67750 6940
rect 67590 5700 67640 6660
rect 67700 5700 67750 6660
rect 67590 5690 67750 5700
rect 67840 7900 68000 7910
rect 67840 6940 67890 7900
rect 67950 6940 68000 7900
rect 67840 6660 68000 6940
rect 67840 5700 67890 6660
rect 67950 5700 68000 6660
rect 67330 4460 67380 5420
rect 67440 4460 67490 5420
rect 67330 4180 67490 4460
rect 67330 3800 67380 4180
rect 67440 3800 67490 4180
rect 67330 3220 67340 3800
rect 67480 3220 67490 3800
rect 67330 3210 67490 3220
rect 67590 5420 67750 5430
rect 67590 4460 67640 5420
rect 67700 4460 67750 5420
rect 67590 4180 67750 4460
rect 67590 3220 67640 4180
rect 67700 3220 67750 4180
rect 67590 3140 67750 3220
rect 67840 5420 68000 5700
rect 67840 4460 67890 5420
rect 67950 4460 68000 5420
rect 67840 4180 68000 4460
rect 67840 3800 67890 4180
rect 67950 3800 68000 4180
rect 67840 3220 67850 3800
rect 67990 3220 68000 3800
rect 67840 3210 68000 3220
rect 68100 7900 68260 7980
rect 68100 6940 68150 7900
rect 68210 6940 68260 7900
rect 68100 6660 68260 6940
rect 68100 5700 68150 6660
rect 68210 5700 68260 6660
rect 68100 5420 68260 5700
rect 68100 4460 68150 5420
rect 68210 4460 68260 5420
rect 68100 4180 68260 4460
rect 68100 3220 68150 4180
rect 68210 3220 68260 4180
rect 68100 3140 68260 3220
rect 68360 7900 68520 7910
rect 68360 6940 68410 7900
rect 68470 6940 68520 7900
rect 68360 6660 68520 6940
rect 68620 7900 68780 7980
rect 68620 6940 68670 7900
rect 68730 6940 68780 7900
rect 68620 6930 68780 6940
rect 68870 7900 69030 7910
rect 68870 6940 68920 7900
rect 68980 6940 69030 7900
rect 68360 5700 68410 6660
rect 68470 5700 68520 6660
rect 68360 5420 68520 5700
rect 68360 4460 68410 5420
rect 68470 4460 68520 5420
rect 68360 4180 68520 4460
rect 68360 3800 68410 4180
rect 68470 3800 68520 4180
rect 68360 3220 68370 3800
rect 68510 3220 68520 3800
rect 68360 3210 68520 3220
rect 68620 6660 68780 6670
rect 68620 5700 68670 6660
rect 68730 5700 68780 6660
rect 68620 5420 68780 5700
rect 68620 4460 68670 5420
rect 68730 4460 68780 5420
rect 68620 4180 68780 4460
rect 68620 3220 68670 4180
rect 68730 3220 68780 4180
rect 68620 3160 68780 3220
rect 68870 6660 69030 6940
rect 68870 5700 68920 6660
rect 68980 5700 69030 6660
rect 68870 5420 69030 5700
rect 69130 7900 69290 7980
rect 69130 6940 69180 7900
rect 69240 6940 69290 7900
rect 69130 6660 69290 6940
rect 69130 5700 69180 6660
rect 69240 5700 69290 6660
rect 69130 5690 69290 5700
rect 69390 7900 69550 7910
rect 69390 6940 69440 7900
rect 69500 6940 69550 7900
rect 69390 6660 69550 6940
rect 69390 5700 69440 6660
rect 69500 5700 69550 6660
rect 68870 4460 68920 5420
rect 68980 4460 69030 5420
rect 68870 4180 69030 4460
rect 68870 3800 68920 4180
rect 68980 3800 69030 4180
rect 68870 3220 68880 3800
rect 69020 3220 69030 3800
rect 68870 3210 69030 3220
rect 69130 5420 69290 5430
rect 69130 4460 69180 5420
rect 69240 4460 69290 5420
rect 69130 4180 69290 4460
rect 69130 3220 69180 4180
rect 69240 3220 69290 4180
rect 60040 2760 67240 3140
rect 67590 2990 68260 3140
rect 68560 2660 68840 3160
rect 69130 3140 69290 3220
rect 69390 5420 69550 5700
rect 69390 4460 69440 5420
rect 69500 4460 69550 5420
rect 69390 4180 69550 4460
rect 69390 3800 69440 4180
rect 69500 3800 69550 4180
rect 69390 3220 69400 3800
rect 69540 3220 69550 3800
rect 69390 3210 69550 3220
rect 69650 7900 69810 7980
rect 69650 6940 69700 7900
rect 69760 6940 69810 7900
rect 69650 6660 69810 6940
rect 69650 5700 69700 6660
rect 69760 5700 69810 6660
rect 69650 5420 69810 5700
rect 69650 4460 69700 5420
rect 69760 4460 69810 5420
rect 69650 4180 69810 4460
rect 69650 3220 69700 4180
rect 69760 3220 69810 4180
rect 69650 3140 69810 3220
rect 69910 7900 70070 7910
rect 69910 6940 69960 7900
rect 70020 6940 70070 7900
rect 69910 6660 70070 6940
rect 70170 7900 70320 7910
rect 70170 6940 70220 7900
rect 70280 6940 70320 7900
rect 70170 6930 70320 6940
rect 70410 7900 70570 7910
rect 70410 6940 70460 7900
rect 70520 6940 70570 7900
rect 69910 5700 69960 6660
rect 70020 5700 70070 6660
rect 69910 5420 70070 5700
rect 69910 4460 69960 5420
rect 70020 4460 70070 5420
rect 69910 4180 70070 4460
rect 69910 3800 69960 4180
rect 70020 3800 70070 4180
rect 69910 3220 69920 3800
rect 70060 3220 70070 3800
rect 69910 3210 70070 3220
rect 70170 6660 70330 6670
rect 70170 5700 70220 6660
rect 70280 5700 70330 6660
rect 70170 5420 70330 5700
rect 70170 4460 70220 5420
rect 70280 4460 70330 5420
rect 70170 4180 70330 4460
rect 70170 3220 70220 4180
rect 70280 3220 70330 4180
rect 70170 3140 70330 3220
rect 70410 6660 70570 6940
rect 70410 5700 70460 6660
rect 70520 5700 70570 6660
rect 70410 5420 70570 5700
rect 70410 4460 70460 5420
rect 70520 4460 70570 5420
rect 70410 4180 70570 4460
rect 70410 3800 70460 4180
rect 70520 3800 70570 4180
rect 70410 3220 70420 3800
rect 70560 3220 70570 3800
rect 70410 3210 70570 3220
rect 70670 7900 70830 8360
rect 71190 8300 71870 8310
rect 71190 8100 71200 8300
rect 71860 8100 71870 8300
rect 71190 7980 71870 8100
rect 70670 6940 70720 7900
rect 70780 6940 70830 7900
rect 70670 6660 70830 6940
rect 70670 5700 70720 6660
rect 70780 5700 70830 6660
rect 70670 5420 70830 5700
rect 70670 4460 70720 5420
rect 70780 4460 70830 5420
rect 70670 4180 70830 4460
rect 70670 3220 70720 4180
rect 70780 3220 70830 4180
rect 70670 3140 70830 3220
rect 70930 7900 71090 7910
rect 70930 6940 70980 7900
rect 71040 6940 71090 7900
rect 70930 6660 71090 6940
rect 70930 5700 70980 6660
rect 71040 5700 71090 6660
rect 70930 5420 71090 5700
rect 71190 7900 71350 7980
rect 71190 6940 71240 7900
rect 71300 6940 71350 7900
rect 71190 6660 71350 6940
rect 71190 5700 71240 6660
rect 71300 5700 71350 6660
rect 71190 5690 71350 5700
rect 71450 7900 71610 7910
rect 71450 6940 71500 7900
rect 71560 6940 71610 7900
rect 71450 6660 71610 6940
rect 71450 5700 71500 6660
rect 71560 5700 71610 6660
rect 70930 4460 70980 5420
rect 71040 4460 71090 5420
rect 70930 4180 71090 4460
rect 70930 3800 70980 4180
rect 71040 3800 71090 4180
rect 70930 3220 70940 3800
rect 71080 3220 71090 3800
rect 70930 3210 71090 3220
rect 71190 5420 71350 5430
rect 71190 4460 71240 5420
rect 71300 4460 71350 5420
rect 71190 4180 71350 4460
rect 71190 3220 71240 4180
rect 71300 3220 71350 4180
rect 71190 3140 71350 3220
rect 71450 5420 71610 5700
rect 71450 4460 71500 5420
rect 71560 4460 71610 5420
rect 71450 4180 71610 4460
rect 71450 3800 71500 4180
rect 71560 3800 71610 4180
rect 71450 3220 71460 3800
rect 71600 3220 71610 3800
rect 71450 3210 71610 3220
rect 71710 7900 71870 7980
rect 72220 7980 74740 8240
rect 71710 6940 71760 7900
rect 71820 6940 71870 7900
rect 71710 6660 71870 6940
rect 71710 5700 71760 6660
rect 71820 5700 71870 6660
rect 71710 5420 71870 5700
rect 71710 4460 71760 5420
rect 71820 4460 71870 5420
rect 71710 4180 71870 4460
rect 71710 3220 71760 4180
rect 71820 3220 71870 4180
rect 71710 3210 71870 3220
rect 71960 7900 72120 7910
rect 71960 6940 72010 7900
rect 72070 6940 72120 7900
rect 71960 6660 72120 6940
rect 71960 5700 72010 6660
rect 72070 5700 72120 6660
rect 71960 5420 72120 5700
rect 71960 4460 72010 5420
rect 72070 4460 72120 5420
rect 71960 4180 72120 4460
rect 71960 3800 72010 4180
rect 72070 3800 72120 4180
rect 71960 3220 71970 3800
rect 72110 3220 72120 3800
rect 71960 3210 72120 3220
rect 72220 7900 72380 7980
rect 72220 6940 72270 7900
rect 72330 6940 72380 7900
rect 72220 6660 72380 6940
rect 72220 5700 72270 6660
rect 72330 5700 72380 6660
rect 72220 5420 72380 5700
rect 72220 4460 72270 5420
rect 72330 4460 72380 5420
rect 72220 4180 72380 4460
rect 72220 3220 72270 4180
rect 72330 3220 72380 4180
rect 69130 2990 69810 3140
rect 59280 2280 68840 2660
rect 70050 2530 70440 3140
rect 70670 2880 71350 3140
rect 72220 3140 72380 3220
rect 72480 7900 72640 7910
rect 72480 6940 72530 7900
rect 72590 6940 72640 7900
rect 72480 6660 72640 6940
rect 72480 5700 72530 6660
rect 72590 5700 72640 6660
rect 72480 5420 72640 5700
rect 72480 4460 72530 5420
rect 72590 4460 72640 5420
rect 72480 4180 72640 4460
rect 72480 3800 72530 4180
rect 72590 3800 72640 4180
rect 72480 3220 72490 3800
rect 72630 3220 72640 3800
rect 72480 3210 72640 3220
rect 72740 7900 72900 7980
rect 72740 6940 72790 7900
rect 72850 6940 72900 7900
rect 72740 6660 72900 6940
rect 72740 5700 72790 6660
rect 72850 5700 72900 6660
rect 72740 5420 72900 5700
rect 72740 4460 72790 5420
rect 72850 4460 72900 5420
rect 72740 4180 72900 4460
rect 72740 3220 72790 4180
rect 72850 3220 72900 4180
rect 72740 3140 72900 3220
rect 73000 7900 73160 7910
rect 73000 6940 73050 7900
rect 73110 6940 73160 7900
rect 73000 6660 73160 6940
rect 73000 5700 73050 6660
rect 73110 5700 73160 6660
rect 73000 5420 73160 5700
rect 73000 4460 73050 5420
rect 73110 4460 73160 5420
rect 73000 4180 73160 4460
rect 73000 3800 73050 4180
rect 73110 3800 73160 4180
rect 73000 3220 73010 3800
rect 73150 3220 73160 3800
rect 73000 3210 73160 3220
rect 73260 7900 73420 7980
rect 73260 6940 73310 7900
rect 73370 6940 73420 7900
rect 73260 6660 73420 6940
rect 73260 5700 73310 6660
rect 73370 5700 73420 6660
rect 73260 5420 73420 5700
rect 73260 4460 73310 5420
rect 73370 4460 73420 5420
rect 73260 4180 73420 4460
rect 73260 3220 73310 4180
rect 73370 3220 73420 4180
rect 73260 3140 73420 3220
rect 73520 7900 73680 7910
rect 73520 6940 73570 7900
rect 73630 6940 73680 7900
rect 73520 6660 73680 6940
rect 73520 5700 73570 6660
rect 73630 5700 73680 6660
rect 73520 5420 73680 5700
rect 73520 4460 73570 5420
rect 73630 4460 73680 5420
rect 73520 4180 73680 4460
rect 74380 4720 74740 7980
rect 74940 6320 75300 8360
rect 81910 8590 82310 8600
rect 81910 8350 81920 8590
rect 82300 8350 82310 8590
rect 81910 8340 82310 8350
rect 74940 5940 75900 6320
rect 83180 6100 83420 8940
rect 90890 8830 91290 9350
rect 84710 8780 85100 8790
rect 84710 8540 84720 8780
rect 85090 8540 85100 8780
rect 84710 7880 85100 8540
rect 86520 8610 91290 8830
rect 84240 7820 84320 7830
rect 84240 6870 84250 7820
rect 84310 6870 84320 7820
rect 83760 6780 84010 6790
rect 83760 6670 83770 6780
rect 84000 6670 84010 6780
rect 83760 6660 84010 6670
rect 84240 6580 84320 6870
rect 83180 6090 83480 6100
rect 83180 5700 83190 6090
rect 83470 5700 83480 6090
rect 83180 5690 83480 5700
rect 84240 5630 84250 6580
rect 84310 5630 84320 6580
rect 84240 5620 84320 5630
rect 84390 7820 84470 7830
rect 84390 6870 84400 7820
rect 84460 6870 84470 7820
rect 84390 6580 84470 6870
rect 84390 5630 84400 6580
rect 84460 5630 84470 6580
rect 84390 5560 84470 5630
rect 84550 7820 84630 7830
rect 84550 6870 84560 7820
rect 84620 6870 84630 7820
rect 84550 6580 84630 6870
rect 84710 7820 84790 7880
rect 84710 6870 84720 7820
rect 84780 6870 84790 7820
rect 84710 6860 84790 6870
rect 84870 7820 84950 7830
rect 84870 6870 84880 7820
rect 84940 6870 84950 7820
rect 84660 6780 84840 6790
rect 84660 6670 84670 6780
rect 84830 6670 84840 6780
rect 84660 6660 84840 6670
rect 84550 5630 84560 6580
rect 84620 5630 84630 6580
rect 84550 5620 84630 5630
rect 84710 6580 84790 6590
rect 84710 5630 84720 6580
rect 84780 5630 84790 6580
rect 84710 5560 84790 5630
rect 84870 6580 84950 6870
rect 84870 5630 84880 6580
rect 84940 5630 84950 6580
rect 84870 5620 84950 5630
rect 85020 7820 85100 7880
rect 85340 7880 86050 7970
rect 85020 6870 85030 7820
rect 85090 6870 85100 7820
rect 85020 6580 85100 6870
rect 85020 5630 85030 6580
rect 85090 5630 85100 6580
rect 85020 5620 85100 5630
rect 85180 7820 85260 7830
rect 85180 6870 85190 7820
rect 85250 6870 85260 7820
rect 85180 6580 85260 6870
rect 85180 5630 85190 6580
rect 85250 5630 85260 6580
rect 85180 5620 85260 5630
rect 85340 7820 85420 7880
rect 85340 6870 85350 7820
rect 85410 6870 85420 7820
rect 85340 6580 85420 6870
rect 85340 5630 85350 6580
rect 85410 5630 85420 6580
rect 84390 5550 84790 5560
rect 84390 5210 84400 5550
rect 84780 5210 84790 5550
rect 85340 5560 85420 5630
rect 85500 7820 85580 7830
rect 85500 6870 85510 7820
rect 85570 6870 85580 7820
rect 85500 6580 85580 6870
rect 85500 5630 85510 6580
rect 85570 5630 85580 6580
rect 85500 5620 85580 5630
rect 85660 7820 85740 7880
rect 85660 6870 85670 7820
rect 85730 6870 85740 7820
rect 85660 6580 85740 6870
rect 85660 5630 85670 6580
rect 85730 5630 85740 6580
rect 85660 5560 85740 5630
rect 85810 7820 85890 7830
rect 85810 6870 85820 7820
rect 85880 6870 85890 7820
rect 85810 6580 85890 6870
rect 85810 5630 85820 6580
rect 85880 5630 85890 6580
rect 85810 5620 85890 5630
rect 85970 7820 86050 7880
rect 85970 6870 85980 7820
rect 86040 6870 86050 7820
rect 85970 6580 86050 6870
rect 85970 5630 85980 6580
rect 86040 5630 86050 6580
rect 85970 5560 86050 5630
rect 86130 7820 86210 7830
rect 86130 6870 86140 7820
rect 86200 6870 86210 7820
rect 86130 6580 86210 6870
rect 86130 5630 86140 6580
rect 86200 5630 86210 6580
rect 86130 5620 86210 5630
rect 85340 5470 86050 5560
rect 84390 5200 84790 5210
rect 86520 4990 86900 8610
rect 84700 4960 85090 4970
rect 74380 4340 76320 4720
rect 73520 3800 73570 4180
rect 73630 3800 73680 4180
rect 73520 3220 73530 3800
rect 73670 3220 73680 3800
rect 73520 3210 73680 3220
rect 72220 2990 73420 3140
rect 79850 2880 80260 4720
rect 84700 4590 84710 4960
rect 85080 4590 85090 4960
rect 84700 4550 85090 4590
rect 69990 2520 70510 2530
rect 69990 2160 70000 2520
rect 70500 2160 70510 2520
rect 70670 2500 80260 2880
rect 84230 4490 84310 4500
rect 84230 3540 84240 4490
rect 84300 3540 84310 4490
rect 84230 3260 84310 3540
rect 84230 2310 84240 3260
rect 84300 2310 84310 3260
rect 84230 2300 84310 2310
rect 84380 4490 84460 4500
rect 84380 3540 84390 4490
rect 84450 3540 84460 4490
rect 84380 3260 84460 3540
rect 84380 2310 84390 3260
rect 84450 2310 84460 3260
rect 69990 2150 70510 2160
rect 84380 2240 84460 2310
rect 84540 4490 84620 4500
rect 84540 3540 84550 4490
rect 84610 3540 84620 4490
rect 84540 3260 84620 3540
rect 84700 4490 84780 4550
rect 84700 3540 84710 4490
rect 84770 3540 84780 4490
rect 84700 3530 84780 3540
rect 84860 4490 84940 4500
rect 84860 3540 84870 4490
rect 84930 3540 84940 4490
rect 84540 2310 84550 3260
rect 84610 2310 84620 3260
rect 84540 2300 84620 2310
rect 84700 3260 84780 3270
rect 84700 2310 84710 3260
rect 84770 2310 84780 3260
rect 84700 2240 84780 2310
rect 84860 3260 84940 3540
rect 84860 2310 84870 3260
rect 84930 2310 84940 3260
rect 84860 2300 84940 2310
rect 85010 4490 85090 4550
rect 85330 4570 86900 4990
rect 85330 4550 86040 4570
rect 85010 3540 85020 4490
rect 85080 3540 85090 4490
rect 85010 3260 85090 3540
rect 85010 2310 85020 3260
rect 85080 2310 85090 3260
rect 85010 2300 85090 2310
rect 85170 4490 85250 4500
rect 85170 3540 85180 4490
rect 85240 3540 85250 4490
rect 85170 3260 85250 3540
rect 85170 2310 85180 3260
rect 85240 2310 85250 3260
rect 85170 2300 85250 2310
rect 85330 4490 85410 4550
rect 85330 3540 85340 4490
rect 85400 3540 85410 4490
rect 85330 3260 85410 3540
rect 85330 2310 85340 3260
rect 85400 2310 85410 3260
rect 84380 2150 84780 2240
rect 85330 2240 85410 2310
rect 85490 4490 85570 4500
rect 85490 3540 85500 4490
rect 85560 3540 85570 4490
rect 85490 3260 85570 3540
rect 85490 2310 85500 3260
rect 85560 2310 85570 3260
rect 85490 2300 85570 2310
rect 85650 4490 85730 4550
rect 85650 3540 85660 4490
rect 85720 3540 85730 4490
rect 85650 3260 85730 3540
rect 85650 2310 85660 3260
rect 85720 2310 85730 3260
rect 85650 2240 85730 2310
rect 85800 4490 85880 4500
rect 85800 3540 85810 4490
rect 85870 3540 85880 4490
rect 85800 3260 85880 3540
rect 85800 2310 85810 3260
rect 85870 2310 85880 3260
rect 85800 2300 85880 2310
rect 85960 4490 86040 4550
rect 85960 3540 85970 4490
rect 86030 3540 86040 4490
rect 85960 3260 86040 3540
rect 85960 2310 85970 3260
rect 86030 2310 86040 3260
rect 85960 2240 86040 2310
rect 86120 4490 86200 4500
rect 86120 3540 86130 4490
rect 86190 3540 86200 4490
rect 86120 3260 86200 3540
rect 86120 2310 86130 3260
rect 86190 2310 86200 3260
rect 93230 3260 93630 3270
rect 93230 2870 93240 3260
rect 93620 2870 93630 3260
rect 93230 2860 93630 2870
rect 86120 2300 86200 2310
rect 85330 2150 86040 2240
rect 50250 2010 50330 2020
rect 41810 1630 54550 1640
rect 41810 1420 54300 1630
rect 54540 1420 54550 1630
rect 41810 1410 54550 1420
rect 52180 1140 52420 1170
rect 52180 1080 54380 1140
rect 51780 1010 52050 1020
rect 51350 920 51600 930
rect 18100 490 20460 840
rect 18100 10 19470 490
rect 20450 10 20460 490
rect 18100 0 20460 10
rect 21840 490 23960 880
rect 21840 10 22970 490
rect 23950 10 23960 490
rect 21840 0 23960 10
rect 25620 490 27820 880
rect 51350 710 51360 920
rect 51590 710 51600 920
rect 51780 850 51790 1010
rect 52040 850 52050 1010
rect 52180 960 52420 1080
rect 54280 1040 54380 1080
rect 52180 900 52190 960
rect 52180 890 52420 900
rect 53390 1030 53630 1040
rect 51780 840 52050 850
rect 53390 840 53400 1030
rect 53620 840 53630 1030
rect 54280 970 54440 1040
rect 53390 830 53630 840
rect 51350 700 51600 710
rect 25620 10 26830 490
rect 27810 10 27820 490
rect 25620 0 27820 10
<< via2 >>
rect 3000 44840 3080 45140
rect 3550 44840 3630 45140
rect 4110 44840 4190 45140
rect 4660 44840 4740 45140
rect 5210 44840 5290 45140
rect 5770 44840 5850 45140
rect 6320 44840 6400 45140
rect 6870 44840 6950 45140
rect 7410 44840 7490 45140
rect 7970 44840 8050 45140
rect 8510 44840 8590 45140
rect 9070 44840 9150 45140
rect 9620 44840 9700 45140
rect 10180 44840 10260 45140
rect 10730 44840 10810 45140
rect 11290 44840 11370 45140
rect 11890 44770 12140 44960
rect 12390 44840 12470 45140
rect 12940 44840 13020 45140
rect 13480 44840 13560 45140
rect 14040 44840 14120 45140
rect 14590 44840 14670 45140
rect 15140 44840 15220 45140
rect 16250 44840 16330 45140
rect 16800 44840 16880 45140
rect 17350 44840 17430 45140
rect 17910 44840 17990 45140
rect 18460 44840 18540 45140
rect 19010 44840 19090 45140
rect 19560 44840 19640 45140
rect 20120 44840 20200 45140
rect 20670 44840 20750 45140
rect 21220 44840 21300 45140
rect 21770 44840 21850 45140
rect 22310 44840 22390 45140
rect 23370 44960 23540 45140
rect 23980 44840 24060 45140
rect 24480 44960 24650 45140
rect 25580 44960 25750 45140
rect 27010 44870 27210 45010
rect 97770 44630 97930 44770
rect 23370 43960 23540 44040
rect 28110 43700 28360 43860
rect 70610 12770 70980 12960
rect 66330 12500 66560 12690
rect 66960 12500 67190 12690
rect 67600 12500 67830 12690
rect 68230 12500 68460 12690
rect 68860 12500 69090 12690
rect 69490 12500 69720 12690
rect 66240 10410 66250 10790
rect 66250 10410 66310 10790
rect 66310 10410 66320 10790
rect 66410 11700 66420 12080
rect 66420 11700 66470 12080
rect 66570 10410 66630 10790
rect 66730 11180 66790 11430
rect 66730 11050 66790 11180
rect 66890 10410 66950 10790
rect 67040 11700 67050 12080
rect 67050 11700 67100 12080
rect 67200 10410 67260 10790
rect 67360 11180 67420 11430
rect 67360 11050 67420 11180
rect 67520 10410 67580 10790
rect 67680 11700 67740 12080
rect 67840 10410 67900 10790
rect 67990 11180 68050 11430
rect 67990 11050 68050 11180
rect 68150 10410 68210 10790
rect 68320 11700 68370 12080
rect 68370 11700 68380 12080
rect 68470 10410 68530 10790
rect 68620 11180 68680 11430
rect 68620 11050 68630 11180
rect 68630 11050 68680 11180
rect 68780 10410 68840 10790
rect 68950 11700 69000 12080
rect 69000 11700 69010 12080
rect 69100 10410 69160 10790
rect 69250 11180 69310 11430
rect 69250 11050 69260 11180
rect 69260 11050 69310 11180
rect 69420 10410 69480 10790
rect 69570 11700 69580 12080
rect 69580 11700 69630 12080
rect 69730 10410 69790 10790
rect 69890 11180 69950 11430
rect 69890 11050 69950 11180
rect 70060 10410 70120 10790
rect 22890 9490 23730 9870
rect 26660 9490 27490 9870
rect 3390 8710 3850 9250
rect 6970 8970 7610 9330
rect 15750 8970 16390 9330
rect 9260 8580 9510 8890
rect 9630 8580 9880 8890
rect 12960 8590 13210 8900
rect 13330 8590 13580 8900
rect 19520 8780 19980 9320
rect 8220 7710 8900 8190
rect 9110 6140 9250 6440
rect 9540 6140 9600 6440
rect 12010 7710 12690 8190
rect 9890 6140 10030 6440
rect 12810 6140 12950 6440
rect 8570 5130 8850 5310
rect 9110 5500 9250 5800
rect 9380 4880 9440 5480
rect 9540 5500 9600 5800
rect 9890 5500 10030 5800
rect 12810 5500 12950 5800
rect 13240 6140 13300 6440
rect 29720 8190 30300 8780
rect 13600 6140 13740 6440
rect 66650 9940 66870 10130
rect 67910 9940 68140 10130
rect 68540 9940 68770 10130
rect 69180 9940 69400 10130
rect 69810 9940 70030 10130
rect 39450 7270 41650 7450
rect 37960 6410 38270 6790
rect 39240 6410 39410 6790
rect 39690 6410 39750 6790
rect 13240 5500 13300 5800
rect 13400 4880 13460 5480
rect 13400 4810 13460 4880
rect 13600 5500 13740 5800
rect 38630 5420 38860 6040
rect 40010 6410 40070 6790
rect 40330 6410 40390 6790
rect 40640 6410 40700 6790
rect 40960 6410 41020 6790
rect 41270 6410 41330 6790
rect 41590 6410 41650 6790
rect 39450 5760 41810 5940
rect 41940 6410 42110 6790
rect 13970 5130 14250 5310
rect 7190 10 8770 390
rect 11350 10 12330 490
rect 15250 10 16230 490
rect 27670 2060 28650 2540
rect 40770 4870 40950 5250
rect 39740 4340 39920 4720
rect 38770 3310 38830 3690
rect 39030 3310 39090 3690
rect 39540 3310 39600 3690
rect 40260 3850 40320 4230
rect 40320 3850 40380 4230
rect 40380 3850 40440 4230
rect 40060 3310 40120 3690
rect 39100 3110 39240 3230
rect 39400 3110 39750 3230
rect 39910 3110 40260 3230
rect 39230 2610 39290 2990
rect 39290 2610 39350 2990
rect 39350 2610 39410 2990
rect 38770 2090 38830 2470
rect 39030 2090 39090 2470
rect 39540 2090 39600 2470
rect 40580 3310 40640 3690
rect 40430 3110 40780 3230
rect 40060 2090 40120 2470
rect 41090 3310 41150 3690
rect 44800 7030 45180 7410
rect 50730 7230 51280 7410
rect 45540 6410 45920 6790
rect 46740 6410 47100 6790
rect 44200 5810 44580 6190
rect 47640 6410 47810 6790
rect 48090 6410 48150 6790
rect 48410 6410 48470 6790
rect 48730 6410 48790 6790
rect 49040 6410 49100 6790
rect 49360 6410 49420 6790
rect 49670 6410 49730 6790
rect 49990 6410 50050 6790
rect 50340 6410 50510 6790
rect 47900 5390 48040 5680
rect 43870 5100 44580 5280
rect 47490 5100 47790 5280
rect 48530 5390 48670 5680
rect 49160 5390 49300 5680
rect 49790 5390 49930 5680
rect 50720 5810 51270 5990
rect 41610 3310 41670 3690
rect 42120 3310 42180 3690
rect 44390 4830 45100 5010
rect 68640 8080 69260 8460
rect 71210 9670 71580 9860
rect 78380 9490 78800 9870
rect 79470 9490 79810 9870
rect 93490 9490 93890 9870
rect 94560 9490 94920 9870
rect 78910 8960 79290 9340
rect 44900 4560 45610 4740
rect 40940 3110 41290 3230
rect 41460 3110 41810 3230
rect 41980 3110 42330 3230
rect 40580 2090 40640 2470
rect 41090 2090 41150 2470
rect 41610 2090 41670 2470
rect 42640 3310 42700 3690
rect 42490 3110 42840 3230
rect 33650 1580 34010 1960
rect 39740 1580 39920 1960
rect 42120 2090 42180 2470
rect 43160 3310 43220 3690
rect 43010 3110 43360 3230
rect 42640 2090 42700 2470
rect 43670 3310 43730 3690
rect 43520 3110 43870 3230
rect 43160 2090 43220 2470
rect 44190 3310 44250 3690
rect 44040 3110 44390 3230
rect 43670 2090 43730 2470
rect 44700 3310 44760 3690
rect 44560 3110 44910 3230
rect 44190 2090 44250 2470
rect 45220 3310 45280 3690
rect 51930 4830 52300 5230
rect 45070 3110 45420 3230
rect 44700 2090 44760 2470
rect 45740 3310 45800 3690
rect 45990 3310 46050 3690
rect 47110 3250 47150 3630
rect 47150 3250 47210 3630
rect 47210 3250 47250 3630
rect 45590 3110 45730 3230
rect 45220 2090 45280 2470
rect 47890 3830 47930 4210
rect 47930 3830 47990 4210
rect 47990 3830 48030 4210
rect 47630 3250 47670 3630
rect 47670 3250 47730 3630
rect 47730 3250 47770 3630
rect 45740 2090 45800 2470
rect 45990 2090 46050 2470
rect 47380 2980 47520 3050
rect 47380 2670 47420 2980
rect 47420 2670 47480 2980
rect 47480 2670 47520 2980
rect 48150 3250 48190 3630
rect 48190 3250 48250 3630
rect 48250 3250 48290 3630
rect 48920 3830 48960 4210
rect 48960 3830 49020 4210
rect 49020 3830 49060 4210
rect 48660 3250 48700 3630
rect 48700 3250 48760 3630
rect 48760 3250 48800 3630
rect 48410 2980 48550 3050
rect 48410 2670 48450 2980
rect 48450 2670 48510 2980
rect 48510 2670 48550 2980
rect 49180 3250 49220 3630
rect 49220 3250 49280 3630
rect 49280 3250 49320 3630
rect 49950 3830 49990 4210
rect 49990 3830 50050 4210
rect 50050 3830 50090 4210
rect 49700 3250 49740 3630
rect 49740 3250 49800 3630
rect 49800 3250 49840 3630
rect 49440 2980 49580 3050
rect 49440 2670 49480 2980
rect 49480 2670 49540 2980
rect 49540 2670 49580 2980
rect 51010 4070 51230 4460
rect 56280 4340 56650 4740
rect 50220 3250 50260 3630
rect 50260 3250 50320 3630
rect 50320 3250 50360 3630
rect 59300 2860 59660 3500
rect 66820 3220 66860 3800
rect 66860 3220 66920 3800
rect 66920 3220 66960 3800
rect 67340 3220 67380 3800
rect 67380 3220 67440 3800
rect 67440 3220 67480 3800
rect 67850 3220 67890 3800
rect 67890 3220 67950 3800
rect 67950 3220 67990 3800
rect 68370 3220 68410 3800
rect 68410 3220 68470 3800
rect 68470 3220 68510 3800
rect 68880 3220 68920 3800
rect 68920 3220 68980 3800
rect 68980 3220 69020 3800
rect 69400 3220 69440 3800
rect 69440 3220 69500 3800
rect 69500 3220 69540 3800
rect 69920 3220 69960 3800
rect 69960 3220 70020 3800
rect 70020 3220 70060 3800
rect 70420 3220 70460 3800
rect 70460 3220 70520 3800
rect 70520 3220 70560 3800
rect 70940 3220 70980 3800
rect 70980 3220 71040 3800
rect 71040 3220 71080 3800
rect 71460 3220 71500 3800
rect 71500 3220 71560 3800
rect 71560 3220 71600 3800
rect 71970 3220 72010 3800
rect 72010 3220 72070 3800
rect 72070 3220 72110 3800
rect 72490 3220 72530 3800
rect 72530 3220 72590 3800
rect 72590 3220 72630 3800
rect 73010 3220 73050 3800
rect 73050 3220 73110 3800
rect 73110 3220 73150 3800
rect 81920 8350 82300 8590
rect 94950 8960 95300 9330
rect 84720 8540 85090 8780
rect 83770 6670 84000 6780
rect 83190 5700 83470 6090
rect 84250 6190 84310 6580
rect 84670 6670 84830 6780
rect 84560 6190 84620 6580
rect 84880 6190 84940 6580
rect 85190 6190 85250 6580
rect 85350 5700 85410 6090
rect 84400 5210 84780 5550
rect 85510 6190 85570 6580
rect 85670 5700 85730 6090
rect 85820 6190 85880 6580
rect 85980 5700 86040 6090
rect 86140 6190 86200 6580
rect 73530 3220 73570 3800
rect 73570 3220 73630 3800
rect 73630 3220 73670 3800
rect 84710 4590 85080 4960
rect 70000 2160 70500 2520
rect 84240 2870 84300 3260
rect 84390 3540 84450 3930
rect 84550 2870 84610 3260
rect 84870 2870 84930 3260
rect 85180 2870 85240 3260
rect 85500 2870 85560 3260
rect 85810 2870 85870 3260
rect 86130 2870 86190 3260
rect 93240 2870 93620 3260
rect 54300 1420 54540 1630
rect 19470 10 20450 490
rect 22970 10 23950 490
rect 51360 710 51590 920
rect 51790 850 52040 1010
rect 53400 840 53620 1030
rect 26830 10 27810 490
<< metal3 >>
rect 2990 45140 3090 45150
rect 2990 44840 3000 45140
rect 3080 44840 3090 45140
rect 2990 44830 3090 44840
rect 3540 45140 3640 45150
rect 3540 44840 3550 45140
rect 3630 44840 3640 45140
rect 3540 44830 3640 44840
rect 4100 45140 4200 45150
rect 4100 44840 4110 45140
rect 4190 44840 4200 45140
rect 4100 44830 4200 44840
rect 4650 45140 4750 45150
rect 4650 44840 4660 45140
rect 4740 44840 4750 45140
rect 4650 44830 4750 44840
rect 5200 45140 5300 45150
rect 5200 44840 5210 45140
rect 5290 44840 5300 45140
rect 5200 44830 5300 44840
rect 5760 45140 5860 45150
rect 5760 44840 5770 45140
rect 5850 44840 5860 45140
rect 5760 44830 5860 44840
rect 6310 45140 6410 45150
rect 6310 44840 6320 45140
rect 6400 44840 6410 45140
rect 6310 44830 6410 44840
rect 6860 45140 6960 45150
rect 6860 44840 6870 45140
rect 6950 44840 6960 45140
rect 6860 44830 6960 44840
rect 7400 45140 7500 45150
rect 7400 44840 7410 45140
rect 7490 44840 7500 45140
rect 7400 44830 7500 44840
rect 7960 45140 8060 45150
rect 7960 44840 7970 45140
rect 8050 44840 8060 45140
rect 7960 44830 8060 44840
rect 8500 45140 8600 45150
rect 8500 44840 8510 45140
rect 8590 44840 8600 45140
rect 8500 44830 8600 44840
rect 9060 45140 9160 45150
rect 9060 44840 9070 45140
rect 9150 44840 9160 45140
rect 9060 44830 9160 44840
rect 9610 45140 9710 45150
rect 9610 44840 9620 45140
rect 9700 44840 9710 45140
rect 9610 44830 9710 44840
rect 10170 45140 10270 45150
rect 10170 44840 10180 45140
rect 10260 44840 10270 45140
rect 10170 44830 10270 44840
rect 10720 45140 10820 45150
rect 10720 44840 10730 45140
rect 10810 44840 10820 45140
rect 10720 44830 10820 44840
rect 11280 45140 11380 45150
rect 11280 44840 11290 45140
rect 11370 44840 11380 45140
rect 12380 45140 12480 45150
rect 11280 44830 11380 44840
rect 11880 44960 12150 44970
rect 11880 44770 11890 44960
rect 12140 44770 12150 44960
rect 12380 44840 12390 45140
rect 12470 44840 12480 45140
rect 12380 44830 12480 44840
rect 12930 45140 13030 45150
rect 12930 44840 12940 45140
rect 13020 44840 13030 45140
rect 12930 44830 13030 44840
rect 13470 45140 13570 45150
rect 13470 44840 13480 45140
rect 13560 44840 13570 45140
rect 13470 44830 13570 44840
rect 14030 45140 14130 45150
rect 14030 44840 14040 45140
rect 14120 44840 14130 45140
rect 14030 44830 14130 44840
rect 14580 45140 14680 45150
rect 14580 44840 14590 45140
rect 14670 44840 14680 45140
rect 14580 44830 14680 44840
rect 15130 45140 15230 45150
rect 15130 44840 15140 45140
rect 15220 44840 15230 45140
rect 15130 44830 15230 44840
rect 16240 45140 16340 45150
rect 16240 44840 16250 45140
rect 16330 44840 16340 45140
rect 16240 44830 16340 44840
rect 16790 45140 16890 45150
rect 16790 44840 16800 45140
rect 16880 44840 16890 45140
rect 16790 44830 16890 44840
rect 17340 45140 17440 45150
rect 17340 44840 17350 45140
rect 17430 44840 17440 45140
rect 17340 44830 17440 44840
rect 17900 45140 18000 45150
rect 17900 44840 17910 45140
rect 17990 44840 18000 45140
rect 17900 44830 18000 44840
rect 18450 45140 18550 45150
rect 18450 44840 18460 45140
rect 18540 44840 18550 45140
rect 18450 44830 18550 44840
rect 19000 45140 19100 45150
rect 19000 44840 19010 45140
rect 19090 44840 19100 45140
rect 19000 44830 19100 44840
rect 19550 45140 19650 45150
rect 19550 44840 19560 45140
rect 19640 44840 19650 45140
rect 19550 44830 19650 44840
rect 20110 45140 20210 45150
rect 20110 44840 20120 45140
rect 20200 44840 20210 45140
rect 20110 44830 20210 44840
rect 20660 45140 20760 45150
rect 20660 44840 20670 45140
rect 20750 44840 20760 45140
rect 20660 44830 20760 44840
rect 21210 45140 21310 45150
rect 21210 44840 21220 45140
rect 21300 44840 21310 45140
rect 21210 44830 21310 44840
rect 21760 45140 21860 45150
rect 21760 44840 21770 45140
rect 21850 44840 21860 45140
rect 21760 44830 21860 44840
rect 22300 45140 22400 45150
rect 22300 44840 22310 45140
rect 22390 44840 22400 45140
rect 23360 45140 23550 45150
rect 23360 44960 23370 45140
rect 23540 44960 23550 45140
rect 23360 44950 23550 44960
rect 23970 45140 24070 45150
rect 22300 44830 22400 44840
rect 23970 44840 23980 45140
rect 24060 44840 24070 45140
rect 24470 45140 24660 45150
rect 24470 44960 24480 45140
rect 24650 44960 24660 45140
rect 24470 44950 24660 44960
rect 25570 45140 25760 45150
rect 25570 44960 25580 45140
rect 25750 44960 25760 45140
rect 25570 44950 25760 44960
rect 27000 45010 27220 45020
rect 27000 44870 27010 45010
rect 27210 44870 27220 45010
rect 27000 44860 27220 44870
rect 23970 44830 24070 44840
rect 11880 44760 12150 44770
rect 15630 44770 15810 44780
rect 15630 44640 15640 44770
rect 97760 44770 97940 44780
rect 97760 44760 97770 44770
rect 15810 44640 97770 44760
rect 15630 44630 97770 44640
rect 97930 44630 97940 44770
rect 15630 44620 97940 44630
rect 170 44420 98260 44430
rect 170 44290 22750 44420
rect 22740 44270 22750 44290
rect 23060 44290 98260 44420
rect 23060 44270 23070 44290
rect 22740 44260 23070 44270
rect 170 44040 98260 44050
rect 170 43960 23370 44040
rect 23540 43960 98260 44040
rect 170 43950 98260 43960
rect 170 43860 98260 43870
rect 170 43750 28110 43860
rect 28100 43700 28110 43750
rect 28360 43750 98260 43860
rect 28360 43700 28370 43750
rect 28100 43690 28370 43700
rect 27310 40380 27550 40390
rect 23220 40370 24260 40380
rect 23450 40190 24260 40370
rect 23220 39990 24260 40190
rect 27310 39760 27320 40380
rect 27540 39990 28140 40380
rect 27540 39760 27550 39990
rect 27310 39560 27550 39760
rect 1880 37800 2280 38660
rect 3340 37960 3940 37970
rect 3340 37800 3350 37960
rect 300 37400 3350 37800
rect 3340 37380 3350 37400
rect 3930 37800 3940 37960
rect 5652 37800 6052 38300
rect 9424 37800 9824 38300
rect 24512 37800 24912 38300
rect 28284 37800 28684 38300
rect 32056 37800 32456 38300
rect 39600 37800 40000 38300
rect 43372 37800 43772 38300
rect 50916 37800 51316 38300
rect 54688 37800 55088 38300
rect 58460 37800 58860 38300
rect 69776 37800 70176 38300
rect 73548 37800 73948 38300
rect 77320 37800 77720 38300
rect 81092 37800 81492 38300
rect 84864 37800 85264 38300
rect 3930 37400 97300 37800
rect 3930 37380 3940 37400
rect 3340 37370 3940 37380
rect 22180 37230 22780 37240
rect 22180 37200 22190 37230
rect 300 36800 13250 37200
rect 13550 36800 17022 37200
rect 17322 36800 20794 37200
rect 21094 36800 22190 37200
rect 22180 36650 22190 36800
rect 22770 37200 22780 37230
rect 22770 36800 35882 37200
rect 36182 37190 47198 37200
rect 36182 36810 41150 37190
rect 41530 36810 47198 37190
rect 36182 36800 47198 36810
rect 47498 36800 62286 37200
rect 62586 36800 66058 37200
rect 66358 36800 88690 37200
rect 88990 36800 92462 37200
rect 92762 36800 96234 37200
rect 96534 36800 97300 37200
rect 22770 36650 22780 36800
rect 22180 36640 22780 36650
rect 300 36610 22100 36618
rect 300 36230 920 36610
rect 1140 36230 4692 36610
rect 4912 36230 8464 36610
rect 8684 36230 12236 36610
rect 12456 36230 16008 36610
rect 16228 36230 19780 36610
rect 20000 36560 22100 36610
rect 22860 36610 97300 36618
rect 22860 36560 23552 36610
rect 20000 36230 23552 36560
rect 23772 36230 27324 36610
rect 27544 36230 31096 36610
rect 31316 36230 34868 36610
rect 35088 36230 38640 36610
rect 38860 36230 42412 36610
rect 42632 36230 46184 36610
rect 46404 36230 49956 36610
rect 50176 36230 53728 36610
rect 53948 36230 57500 36610
rect 57720 36230 61272 36610
rect 61492 36230 65044 36610
rect 65264 36230 68816 36610
rect 69036 36230 72588 36610
rect 72808 36230 76360 36610
rect 76580 36230 80132 36610
rect 80352 36230 83904 36610
rect 84124 36230 87676 36610
rect 87896 36230 91448 36610
rect 91668 36230 95220 36610
rect 95440 36230 97300 36610
rect 300 36220 97300 36230
rect 27310 35758 27550 35768
rect 23220 35748 24260 35758
rect 23450 35568 24260 35748
rect 23220 35368 24260 35568
rect 27310 35138 27320 35758
rect 27540 35368 28140 35758
rect 27540 35138 27550 35368
rect 27310 34938 27550 35138
rect 1880 33178 2280 34038
rect 5652 33178 6052 33678
rect 7110 33300 7710 33310
rect 7110 33178 7120 33300
rect 300 32778 7120 33178
rect 7110 32720 7120 32778
rect 7700 33178 7710 33300
rect 9424 33178 9824 33678
rect 24512 33178 24912 33678
rect 28284 33178 28684 33678
rect 32056 33178 32456 33678
rect 39600 33178 40000 33678
rect 43372 33178 43772 33678
rect 50916 33178 51316 33678
rect 54688 33178 55088 33678
rect 58460 33178 58860 33678
rect 69776 33178 70176 33678
rect 73548 33178 73948 33678
rect 77320 33178 77720 33678
rect 81092 33178 81492 33678
rect 84864 33178 85264 33678
rect 7700 32778 97300 33178
rect 7700 32720 7710 32778
rect 7110 32710 7710 32720
rect 25970 32610 26570 32620
rect 25970 32578 25980 32610
rect 300 32178 13250 32578
rect 13550 32178 17022 32578
rect 17322 32178 20794 32578
rect 21094 32178 25980 32578
rect 25970 32030 25980 32178
rect 26560 32578 26570 32610
rect 26560 32178 35882 32578
rect 36182 32178 47198 32578
rect 47498 32570 62286 32578
rect 47498 32190 48700 32570
rect 49070 32190 62286 32570
rect 47498 32178 62286 32190
rect 62586 32178 66058 32578
rect 66358 32178 88690 32578
rect 88990 32178 92462 32578
rect 92762 32178 96234 32578
rect 96534 32178 97300 32578
rect 26560 32030 26570 32178
rect 25970 32020 26570 32030
rect 27310 31136 27550 31146
rect 23220 31126 24260 31136
rect 23450 30946 24260 31126
rect 23220 30746 24260 30946
rect 27310 30516 27320 31136
rect 27540 30746 28140 31136
rect 27540 30516 27550 30746
rect 27310 30316 27550 30516
rect 1880 28556 2280 29416
rect 5652 28556 6052 29056
rect 9424 28556 9824 29056
rect 10890 28680 11490 28690
rect 10890 28556 10900 28680
rect 300 28156 10900 28556
rect 10890 28100 10900 28156
rect 11480 28556 11490 28680
rect 24512 28556 24912 29056
rect 28284 28556 28684 29056
rect 32056 28556 32456 29056
rect 39600 28556 40000 29056
rect 43372 28556 43772 29056
rect 50916 28556 51316 29056
rect 54688 28556 55088 29056
rect 58460 28556 58860 29056
rect 69776 28556 70176 29056
rect 73548 28556 73948 29056
rect 77320 28556 77720 29056
rect 81092 28556 81492 29056
rect 84864 28556 85264 29056
rect 11480 28156 97300 28556
rect 11480 28100 11490 28156
rect 10890 28090 11490 28100
rect 29720 28020 30320 28030
rect 29720 27956 29730 28020
rect 300 27556 13250 27956
rect 13550 27556 17022 27956
rect 17322 27556 20794 27956
rect 21094 27556 29730 27956
rect 29720 27440 29730 27556
rect 30310 27956 30320 28020
rect 30310 27556 35882 27956
rect 36182 27556 47198 27956
rect 47498 27940 62286 27956
rect 47498 27570 56240 27940
rect 56620 27570 62286 27940
rect 47498 27556 62286 27570
rect 62586 27556 66058 27956
rect 66358 27556 88690 27956
rect 88990 27556 92462 27956
rect 92762 27556 96234 27956
rect 96534 27556 97300 27956
rect 30310 27440 30320 27556
rect 29720 27430 30320 27440
rect 27310 26514 27550 26524
rect 23220 26504 24260 26514
rect 23450 26324 24260 26504
rect 23220 26124 24260 26324
rect 27310 25894 27320 26514
rect 27540 26124 28140 26514
rect 27540 25894 27550 26124
rect 27310 25694 27550 25894
rect 1880 23934 2280 24794
rect 5652 23934 6052 24434
rect 9424 23934 9824 24434
rect 14660 24060 15260 24070
rect 14660 23934 14670 24060
rect 300 23534 14670 23934
rect 14660 23480 14670 23534
rect 15250 23934 15260 24060
rect 24512 23934 24912 24434
rect 28284 23934 28684 24434
rect 32056 23934 32456 24434
rect 39600 23934 40000 24434
rect 54688 23934 55088 24434
rect 58460 23934 58860 24434
rect 73548 23934 73948 24434
rect 77320 23934 77720 24434
rect 81092 23934 81492 24434
rect 84864 23934 85264 24434
rect 90130 24150 90660 24160
rect 90130 23934 90140 24150
rect 15250 23534 90140 23934
rect 15250 23480 15260 23534
rect 14660 23470 15260 23480
rect 90130 23470 90140 23534
rect 90650 23934 90660 24150
rect 90650 23534 97300 23934
rect 90650 23470 90660 23534
rect 90130 23460 90660 23470
rect 75120 23370 75520 23380
rect 75120 23334 75130 23370
rect 300 22934 13250 23334
rect 13550 22934 17022 23334
rect 17322 22934 20794 23334
rect 21094 22934 35882 23334
rect 36182 22934 47198 23334
rect 47498 22934 62286 23334
rect 62586 22934 66058 23334
rect 66358 22934 75130 23334
rect 39460 22730 43426 22740
rect 39460 22350 41150 22730
rect 41530 22350 43426 22730
rect 39460 22340 43426 22350
rect 43726 22340 50970 22740
rect 51270 22340 69830 22740
rect 70130 22340 71780 22740
rect 75120 22390 75130 22934
rect 75520 22934 88690 23334
rect 88990 22934 92462 23334
rect 92762 22934 96234 23334
rect 96534 22934 97300 23334
rect 75120 22380 75520 22390
rect 27310 21892 27550 21902
rect 23220 21882 24260 21892
rect 23450 21702 24260 21882
rect 23220 21502 24260 21702
rect 27310 21272 27320 21892
rect 27540 21502 28140 21892
rect 27540 21272 27550 21502
rect 27310 21072 27550 21272
rect 1880 19312 2280 20172
rect 5652 19312 6052 19812
rect 9424 19312 9824 19812
rect 18420 19440 19020 19450
rect 18420 19312 18430 19440
rect 300 18912 18430 19312
rect 18420 18860 18430 18912
rect 19010 19312 19020 19440
rect 24512 19312 24912 19812
rect 28284 19312 28684 19812
rect 32056 19312 32456 19812
rect 39600 19312 40000 19812
rect 54688 19312 55088 19812
rect 58460 19312 58860 19812
rect 73548 19312 73948 19812
rect 77320 19312 77720 19812
rect 81092 19312 81492 19812
rect 84864 19312 85264 19812
rect 93900 19520 94430 19530
rect 93900 19312 93910 19520
rect 19010 18912 93910 19312
rect 19010 18860 19020 18912
rect 18420 18850 19020 18860
rect 93900 18840 93910 18912
rect 94420 19312 94430 19520
rect 94420 18912 97300 19312
rect 94420 18840 94430 18912
rect 93900 18830 94430 18840
rect 78900 18740 79300 18750
rect 78900 18712 78910 18740
rect 300 18312 13250 18712
rect 13550 18312 17022 18712
rect 17322 18312 20794 18712
rect 21094 18312 35882 18712
rect 36182 18312 47198 18712
rect 47498 18312 62286 18712
rect 62586 18312 66058 18712
rect 66358 18312 78910 18712
rect 39460 17718 43426 18118
rect 43726 18110 50970 18118
rect 43726 17730 48700 18110
rect 49070 17730 50970 18110
rect 43726 17718 50970 17730
rect 51270 17718 69830 18118
rect 70130 17718 71780 18118
rect 78900 17760 78910 18312
rect 79290 18712 79300 18740
rect 79290 18312 88690 18712
rect 88990 18312 92462 18712
rect 92762 18312 96234 18712
rect 96534 18312 97300 18712
rect 79290 17760 79300 18312
rect 78900 17750 79300 17760
rect 27310 17270 27550 17280
rect 23220 17260 24490 17270
rect 23450 17080 24490 17260
rect 23220 16880 24490 17080
rect 27310 16650 27320 17270
rect 27540 16880 28140 17270
rect 27540 16650 27550 16880
rect 27310 16450 27550 16650
rect 1880 14690 2280 15550
rect 5652 14690 6052 15190
rect 9424 14690 9824 15190
rect 24512 14690 24912 15190
rect 28284 14690 28684 15190
rect 32056 14690 32456 15190
rect 39600 14690 40000 15190
rect 54688 14690 55088 15190
rect 58460 14690 58860 15190
rect 73548 14690 73948 15190
rect 77320 14690 77720 15190
rect 81092 14690 81492 15190
rect 84864 14690 85264 15190
rect 300 14680 98160 14690
rect 300 14290 97770 14680
rect 82670 14090 83070 14100
rect 300 13690 13250 14090
rect 13550 13690 17022 14090
rect 17322 13690 20794 14090
rect 21094 13690 35882 14090
rect 36182 13690 47198 14090
rect 47498 13690 62286 14090
rect 62586 13690 66058 14090
rect 66358 13690 82680 14090
rect 39460 13096 43426 13496
rect 43726 13096 50970 13496
rect 51270 13480 69830 13496
rect 51270 13110 56240 13480
rect 56610 13110 69830 13480
rect 51270 13096 69830 13110
rect 70130 13096 71780 13496
rect 82670 13110 82680 13690
rect 83060 13690 88690 14090
rect 88990 13690 92462 14090
rect 92762 13690 96234 14090
rect 96534 13690 97300 14090
rect 97760 13700 97770 14290
rect 98150 13700 98160 14680
rect 97760 13690 98160 13700
rect 83060 13110 83070 13690
rect 82670 13100 83070 13110
rect 70600 12960 70990 12970
rect 25260 12840 25860 12850
rect 25260 12260 25270 12840
rect 25850 12260 25860 12840
rect 25260 12250 25860 12260
rect 29080 12840 29680 12850
rect 29080 12260 29090 12840
rect 29670 12260 29680 12840
rect 70600 12770 70610 12960
rect 70980 12770 70990 12960
rect 70600 12760 70990 12770
rect 66230 12690 71590 12700
rect 66230 12500 66330 12690
rect 66560 12500 66960 12690
rect 67190 12500 67600 12690
rect 67830 12500 68230 12690
rect 68460 12500 68860 12690
rect 69090 12500 69490 12690
rect 69720 12500 71210 12690
rect 71580 12500 71590 12690
rect 66230 12490 71590 12500
rect 29080 12250 29680 12260
rect 66230 12080 71810 12090
rect 66230 11700 66410 12080
rect 66470 11700 67040 12080
rect 67100 11700 67680 12080
rect 67740 11700 68320 12080
rect 68380 11700 68950 12080
rect 69010 11700 69570 12080
rect 69630 11700 71810 12080
rect 66230 11690 71810 11700
rect 66230 11430 70150 11440
rect 66230 11050 66730 11430
rect 66790 11050 66840 11430
rect 67210 11050 67360 11430
rect 67420 11050 67990 11430
rect 68050 11050 68620 11430
rect 68680 11050 69250 11430
rect 69310 11050 69890 11430
rect 69950 11050 70150 11430
rect 66230 11040 70150 11050
rect 3110 10330 3380 10950
rect 4020 10330 4290 10950
rect 3110 10120 4290 10330
rect 18190 10330 18460 10550
rect 19110 10330 19380 10550
rect 66230 10790 70150 10800
rect 66230 10410 66240 10790
rect 66320 10410 66570 10790
rect 66630 10410 66890 10790
rect 66950 10410 67200 10790
rect 67260 10410 67520 10790
rect 67580 10410 67840 10790
rect 67900 10410 68150 10790
rect 68210 10410 68470 10790
rect 68530 10410 68780 10790
rect 68840 10410 69100 10790
rect 69160 10410 69420 10790
rect 69480 10410 69730 10790
rect 69790 10410 70060 10790
rect 70120 10410 70150 10790
rect 66230 10400 70150 10410
rect 71440 10420 71810 11690
rect 71440 10410 74760 10420
rect 18190 10120 19380 10330
rect 66230 10130 70990 10140
rect 26080 10060 26480 10070
rect 22320 10030 22720 10040
rect 22320 9340 22330 10030
rect 22710 9880 22720 10030
rect 22710 9870 23740 9880
rect 22710 9490 22890 9870
rect 23730 9490 23740 9870
rect 22710 9480 23740 9490
rect 22710 9340 22720 9480
rect 26080 9370 26090 10060
rect 26470 9880 26480 10060
rect 66230 9940 66650 10130
rect 66870 9940 67910 10130
rect 68140 9940 68540 10130
rect 68770 9940 69180 10130
rect 69400 9940 69810 10130
rect 70030 9940 70610 10130
rect 70980 9940 70990 10130
rect 71440 10020 74380 10410
rect 74750 10020 74760 10410
rect 71440 10010 74760 10020
rect 66230 9930 70990 9940
rect 26470 9870 27500 9880
rect 78370 9870 79820 9880
rect 26470 9490 26660 9870
rect 27490 9490 27500 9870
rect 71200 9860 71590 9870
rect 71200 9670 71210 9860
rect 71580 9670 71590 9860
rect 71200 9660 71590 9670
rect 26470 9480 27500 9490
rect 78370 9490 78380 9870
rect 78800 9490 79470 9870
rect 79810 9490 79820 9870
rect 78370 9480 79820 9490
rect 93480 9870 94930 9880
rect 93480 9490 93490 9870
rect 93890 9490 94560 9870
rect 94920 9490 94930 9870
rect 93480 9480 94930 9490
rect 26470 9370 26480 9480
rect 26080 9360 26480 9370
rect 6960 9330 7620 9340
rect 3380 9250 3860 9260
rect 3380 8710 3390 9250
rect 3850 8900 3860 9250
rect 6960 8970 6970 9330
rect 7610 9180 7620 9330
rect 15740 9330 16400 9340
rect 22320 9330 22720 9340
rect 78890 9340 85110 9350
rect 15740 9190 15750 9330
rect 7610 8980 9890 9180
rect 7610 8970 7620 8980
rect 6960 8960 7620 8970
rect 3850 8890 9520 8900
rect 3850 8710 9260 8890
rect 3380 8700 9260 8710
rect 9250 8580 9260 8700
rect 9510 8580 9520 8890
rect 9250 8570 9520 8580
rect 9620 8890 9890 8980
rect 9620 8580 9630 8890
rect 9880 8580 9890 8890
rect 12950 8990 15750 9190
rect 12950 8900 13220 8990
rect 15740 8970 15750 8990
rect 16390 8970 16400 9330
rect 15740 8960 16400 8970
rect 19510 9320 19990 9330
rect 12950 8590 12960 8900
rect 13210 8590 13220 8900
rect 12950 8580 13220 8590
rect 13320 8900 13590 8910
rect 19510 8900 19520 9320
rect 13320 8590 13330 8900
rect 13580 8780 19520 8900
rect 19980 8780 19990 9320
rect 78890 8960 78910 9340
rect 79290 8960 85110 9340
rect 78890 8950 85110 8960
rect 86520 9340 95320 9350
rect 86520 8960 86530 9340
rect 86880 9330 95320 9340
rect 86880 8960 94950 9330
rect 95300 8960 95320 9330
rect 86520 8950 95320 8960
rect 13580 8700 19990 8780
rect 29710 8780 30310 8790
rect 13580 8590 13590 8700
rect 13320 8580 13590 8590
rect 9620 8570 9890 8580
rect 8200 8190 8920 8200
rect 8200 7710 8220 8190
rect 8900 7710 8920 8190
rect 8200 7700 8920 7710
rect 12000 8190 12700 8200
rect 12000 7710 12010 8190
rect 12690 7710 12700 8190
rect 29710 8190 29720 8780
rect 30300 8190 30310 8780
rect 84710 8780 85110 8950
rect 81910 8590 82310 8600
rect 29710 8180 30310 8190
rect 63040 8160 63060 8480
rect 63440 8460 69280 8480
rect 63440 8160 68640 8460
rect 68620 8080 68640 8160
rect 69260 8080 69280 8460
rect 81910 8350 81920 8590
rect 82300 8350 82310 8590
rect 84710 8540 84720 8780
rect 85090 8540 85110 8780
rect 84710 8530 85110 8540
rect 81910 8340 82310 8350
rect 68620 8060 69280 8080
rect 47960 7860 47980 8050
rect 12000 7700 12700 7710
rect 43310 7670 47980 7860
rect 48350 7670 48370 8050
rect 43310 7660 48370 7670
rect 43310 7460 43530 7660
rect 52330 7610 52730 7620
rect 39440 7450 43530 7460
rect 39440 7270 39450 7450
rect 41650 7270 43530 7450
rect 39440 7260 43530 7270
rect 44790 7410 45190 7460
rect 52330 7420 52340 7610
rect 44790 7030 44800 7410
rect 45180 7030 45190 7410
rect 50720 7410 52340 7420
rect 50720 7230 50730 7410
rect 51280 7230 52340 7410
rect 52720 7230 52730 7610
rect 50720 7220 52730 7230
rect 44790 7020 45190 7030
rect 37950 6790 45930 6800
rect 9100 6440 9260 6450
rect 9100 6140 9110 6440
rect 9250 6350 9260 6440
rect 9530 6440 9610 6450
rect 9530 6350 9540 6440
rect 9250 6150 9540 6350
rect 9250 6140 9260 6150
rect 9100 6130 9260 6140
rect 9530 6140 9540 6150
rect 9600 6350 9610 6440
rect 9880 6440 10040 6450
rect 9880 6350 9890 6440
rect 9600 6150 9890 6350
rect 9600 6140 9610 6150
rect 9530 6130 9610 6140
rect 9880 6140 9890 6150
rect 10030 6350 10040 6440
rect 12800 6440 12960 6450
rect 10240 6350 10650 6360
rect 10030 6150 10250 6350
rect 10030 6140 10040 6150
rect 9880 6130 10040 6140
rect 9100 5800 9260 5810
rect 9100 5500 9110 5800
rect 9250 5790 9260 5800
rect 9530 5800 9610 5810
rect 9530 5790 9540 5800
rect 9250 5590 9540 5790
rect 9250 5500 9260 5590
rect 9100 5490 9260 5500
rect 9530 5500 9540 5590
rect 9600 5790 9610 5800
rect 9880 5800 10040 5810
rect 9880 5790 9890 5800
rect 9600 5590 9890 5790
rect 9600 5500 9610 5590
rect 9530 5490 9610 5500
rect 9880 5500 9890 5590
rect 10030 5790 10040 5800
rect 10240 5790 10250 6150
rect 10030 5590 10250 5790
rect 10640 5590 10650 6350
rect 12800 6140 12810 6440
rect 12950 6350 12960 6440
rect 13230 6440 13310 6450
rect 13230 6350 13240 6440
rect 12950 6150 13240 6350
rect 12950 6140 12960 6150
rect 12800 6130 12960 6140
rect 13230 6140 13240 6150
rect 13300 6350 13310 6440
rect 13590 6440 13750 6450
rect 13590 6350 13600 6440
rect 13300 6150 13600 6350
rect 13300 6140 13310 6150
rect 13230 6130 13310 6140
rect 13590 6140 13600 6150
rect 13740 6350 13750 6440
rect 37950 6410 37960 6790
rect 38270 6410 39240 6790
rect 39410 6410 39690 6790
rect 39750 6410 40010 6790
rect 40070 6410 40330 6790
rect 40390 6410 40640 6790
rect 40700 6410 40960 6790
rect 41020 6410 41270 6790
rect 41330 6410 41590 6790
rect 41650 6410 41940 6790
rect 42110 6410 45540 6790
rect 45920 6410 45930 6790
rect 37950 6400 45930 6410
rect 46170 6790 47110 6800
rect 46170 6410 46180 6790
rect 46430 6410 46740 6790
rect 47100 6410 47110 6790
rect 46170 6400 47110 6410
rect 47630 6790 50530 6800
rect 47630 6410 47640 6790
rect 47810 6410 48090 6790
rect 48150 6410 48410 6790
rect 48470 6410 48730 6790
rect 48790 6410 49040 6790
rect 49100 6410 49360 6790
rect 49420 6410 49670 6790
rect 49730 6410 49990 6790
rect 50050 6410 50340 6790
rect 50510 6410 50530 6790
rect 83760 6780 84860 6790
rect 83760 6670 83770 6780
rect 84000 6670 84670 6780
rect 84830 6670 84860 6780
rect 83760 6660 84860 6670
rect 47630 6400 50530 6410
rect 84230 6580 86220 6590
rect 14010 6350 14420 6360
rect 13740 6150 14020 6350
rect 13740 6140 13750 6150
rect 13590 6130 13750 6140
rect 10030 5500 10040 5590
rect 10240 5580 10650 5590
rect 12800 5800 12960 5810
rect 9880 5490 10040 5500
rect 12800 5500 12810 5800
rect 12950 5790 12960 5800
rect 13230 5800 13310 5810
rect 13230 5790 13240 5800
rect 12950 5590 13240 5790
rect 12950 5500 12960 5590
rect 12800 5490 12960 5500
rect 13230 5500 13240 5590
rect 13300 5790 13310 5800
rect 13590 5800 13750 5810
rect 13590 5790 13600 5800
rect 13300 5590 13600 5790
rect 13300 5500 13310 5590
rect 13230 5490 13310 5500
rect 13590 5500 13600 5590
rect 13740 5790 13750 5800
rect 14010 5790 14020 6150
rect 13740 5590 14020 5790
rect 14410 5590 14420 6350
rect 44190 6190 44590 6200
rect 38620 6040 38870 6050
rect 13740 5500 13750 5590
rect 14010 5580 14420 5590
rect 13590 5490 13750 5500
rect 9370 5480 9450 5490
rect 6460 5310 8860 5320
rect 6460 5130 6480 5310
rect 6860 5130 8570 5310
rect 8850 5130 8860 5310
rect 6460 5120 8860 5130
rect 9370 5000 9380 5480
rect 2700 4990 9380 5000
rect 2700 4810 2710 4990
rect 3090 4880 9380 4990
rect 9440 4880 9450 5480
rect 3090 4810 9450 4880
rect 2700 4800 9450 4810
rect 13390 5480 13470 5490
rect 13390 4810 13400 5480
rect 13460 5000 13470 5480
rect 38620 5420 38630 6040
rect 38860 5420 38870 6040
rect 39440 5940 41820 5950
rect 39440 5760 39450 5940
rect 41810 5760 41820 5940
rect 44190 5810 44200 6190
rect 44580 5810 44590 6190
rect 51730 6190 52130 6200
rect 51730 6000 51740 6190
rect 44190 5800 44590 5810
rect 50710 5990 51740 6000
rect 50710 5810 50720 5990
rect 51270 5810 51740 5990
rect 52120 5810 52130 6190
rect 84230 6190 84250 6580
rect 84310 6190 84560 6580
rect 84620 6190 84880 6580
rect 84940 6190 85190 6580
rect 85250 6190 85510 6580
rect 85570 6190 85690 6580
rect 86070 6190 86140 6580
rect 86200 6190 86220 6580
rect 84230 6180 86220 6190
rect 83180 6090 86090 6100
rect 50710 5800 52130 5810
rect 39440 5750 40430 5760
rect 40420 5560 40430 5750
rect 40810 5750 41820 5760
rect 40810 5560 40820 5750
rect 55510 5740 55910 5750
rect 55510 5690 55520 5740
rect 40420 5550 40820 5560
rect 47860 5680 55520 5690
rect 38620 5410 38870 5420
rect 47860 5390 47900 5680
rect 48040 5390 48530 5680
rect 48670 5390 49160 5680
rect 49300 5390 49790 5680
rect 49930 5390 50660 5680
rect 50880 5390 55520 5680
rect 55900 5390 55910 5740
rect 83180 5700 83190 6090
rect 83470 5700 85350 6090
rect 85410 5700 85670 6090
rect 85730 5700 85980 6090
rect 86040 5700 86090 6090
rect 83180 5690 86090 5700
rect 47860 5380 55910 5390
rect 78140 5550 84790 5560
rect 13960 5310 17790 5320
rect 13960 5130 13970 5310
rect 14250 5130 17790 5310
rect 13960 5120 17790 5130
rect 18180 5120 18200 5320
rect 43860 5280 47800 5290
rect 37410 5250 40960 5260
rect 13460 4810 21570 5000
rect 13390 4800 21570 4810
rect 21950 4800 21960 5000
rect 37410 4870 37420 5250
rect 37790 4870 40770 5250
rect 40950 4870 40960 5250
rect 43860 5100 43870 5280
rect 44580 5100 47490 5280
rect 47790 5100 47800 5280
rect 43860 5090 47800 5100
rect 51920 5230 52310 5240
rect 51920 5020 51930 5230
rect 37410 4860 40960 4870
rect 44380 5010 51930 5020
rect 44380 4830 44390 5010
rect 45100 4830 51930 5010
rect 52300 4830 52310 5230
rect 78140 5210 78150 5550
rect 78530 5210 84400 5550
rect 84780 5210 84790 5550
rect 78140 5200 84790 5210
rect 44380 4820 52310 4830
rect 84700 4960 86890 4970
rect 44890 4740 56660 4750
rect 36640 4720 39930 4730
rect 36640 4340 36650 4720
rect 37040 4340 39740 4720
rect 39920 4340 39930 4720
rect 44890 4560 44900 4740
rect 45610 4560 56280 4740
rect 44890 4550 56280 4560
rect 36640 4330 39930 4340
rect 51000 4460 51240 4470
rect 33640 4230 40450 4240
rect 24050 3950 25050 3960
rect 24050 3900 24060 3950
rect 1350 3890 24060 3900
rect 1350 3500 3150 3890
rect 3140 3410 3150 3500
rect 3860 3500 24060 3890
rect 3860 3410 4140 3500
rect 24050 3470 24060 3500
rect 25040 3900 25050 3950
rect 25040 3500 30050 3900
rect 33640 3850 33650 4230
rect 34020 3850 40260 4230
rect 40440 3850 40450 4230
rect 33640 3840 40450 3850
rect 47140 4210 50890 4220
rect 47140 3830 47890 4210
rect 48030 3830 48920 4210
rect 49060 3830 49950 4210
rect 50090 3830 50660 4210
rect 50880 3830 50890 4210
rect 51000 4070 51010 4460
rect 51230 4070 51240 4460
rect 56270 4340 56280 4550
rect 56650 4340 56660 4740
rect 84700 4590 84710 4960
rect 85080 4590 86530 4960
rect 86880 4590 86890 4960
rect 84700 4580 86890 4590
rect 56270 4330 56660 4340
rect 51000 4060 51240 4070
rect 84220 4040 86210 4450
rect 47140 3820 50890 3830
rect 84220 3930 97400 3940
rect 65030 3800 73680 3810
rect 38220 3690 46060 3700
rect 25040 3470 25050 3500
rect 24050 3460 25050 3470
rect 3140 3400 4140 3410
rect 38220 3310 38310 3690
rect 38540 3310 38770 3690
rect 38830 3310 39030 3690
rect 39090 3310 39540 3690
rect 39600 3310 40060 3690
rect 40120 3310 40580 3690
rect 40640 3310 41090 3690
rect 41150 3310 41610 3690
rect 41670 3310 42120 3690
rect 42180 3310 42640 3690
rect 42700 3310 43160 3690
rect 43220 3310 43670 3690
rect 43730 3310 44190 3690
rect 44250 3310 44700 3690
rect 44760 3310 45220 3690
rect 45280 3310 45740 3690
rect 45800 3310 45990 3690
rect 46050 3310 46060 3690
rect 38220 3300 46060 3310
rect 46170 3630 50370 3640
rect 6900 3250 7900 3260
rect 46170 3250 46180 3630
rect 46610 3250 47110 3630
rect 47250 3250 47630 3630
rect 47770 3250 48150 3630
rect 48290 3250 48660 3630
rect 48800 3250 49180 3630
rect 49320 3250 49700 3630
rect 49840 3250 50220 3630
rect 50360 3250 50370 3630
rect 6900 3200 6910 3250
rect 1350 2800 6910 3200
rect 6900 2770 6910 2800
rect 7620 3200 7900 3250
rect 20430 3240 21430 3250
rect 20430 3200 20440 3240
rect 7620 2800 20440 3200
rect 7620 2770 7900 2800
rect 6900 2760 7900 2770
rect 20430 2760 20440 2800
rect 21420 3200 21430 3240
rect 28860 3240 29860 3250
rect 46170 3240 50370 3250
rect 59280 3500 59680 3520
rect 28860 3200 28870 3240
rect 21420 2800 28870 3200
rect 21420 2760 21430 2800
rect 20430 2750 21430 2760
rect 28860 2760 28870 2800
rect 29850 3200 29860 3240
rect 32640 3230 45750 3240
rect 29850 2800 30050 3200
rect 32640 3110 39100 3230
rect 39240 3110 39400 3230
rect 39750 3110 39910 3230
rect 40260 3110 40430 3230
rect 40780 3110 40940 3230
rect 41290 3110 41460 3230
rect 41810 3110 41980 3230
rect 42330 3110 42490 3230
rect 42840 3110 43010 3230
rect 43360 3110 43520 3230
rect 43870 3110 44040 3230
rect 44390 3110 44560 3230
rect 44910 3110 45070 3230
rect 45420 3110 45590 3230
rect 45730 3110 45750 3230
rect 32640 3100 45750 3110
rect 47140 3050 54810 3060
rect 32870 2990 39420 3000
rect 29850 2760 29860 2800
rect 28860 2750 29860 2760
rect 32870 2610 32880 2990
rect 33270 2610 39230 2990
rect 39410 2610 39420 2990
rect 47140 2670 47380 3050
rect 47520 2670 48410 3050
rect 48550 2670 49440 3050
rect 49580 2670 54810 3050
rect 59280 2860 59300 3500
rect 59660 2860 59680 3500
rect 65030 3220 65040 3800
rect 65480 3220 66820 3800
rect 66960 3220 67340 3800
rect 67480 3220 67850 3800
rect 67990 3220 68370 3800
rect 68510 3220 68880 3800
rect 69020 3220 69400 3800
rect 69540 3220 69920 3800
rect 70060 3220 70420 3800
rect 70560 3220 70940 3800
rect 71080 3220 71460 3800
rect 71600 3220 71970 3800
rect 72110 3220 72490 3800
rect 72630 3220 73010 3800
rect 73150 3220 73530 3800
rect 73670 3220 73680 3800
rect 84220 3540 84390 3930
rect 84450 3540 97010 3930
rect 84220 3530 97010 3540
rect 97390 3530 97400 3930
rect 97000 3520 97400 3530
rect 65030 3210 73680 3220
rect 84220 3260 89860 3270
rect 84220 2870 84240 3260
rect 84300 2870 84550 3260
rect 84610 2870 84870 3260
rect 84930 2870 85180 3260
rect 85240 2870 85500 3260
rect 85560 2870 85810 3260
rect 85870 2870 86130 3260
rect 86190 2870 89470 3260
rect 89840 2870 89860 3260
rect 84220 2860 89860 2870
rect 93230 3260 93630 3270
rect 93230 2870 93240 3260
rect 93620 2870 93630 3260
rect 93230 2860 93630 2870
rect 59280 2840 59680 2860
rect 47140 2660 54810 2670
rect 32870 2600 39420 2610
rect 10700 2550 11700 2560
rect 10700 2500 10710 2550
rect 1350 2100 10710 2500
rect 10700 2070 10710 2100
rect 11420 2500 11700 2550
rect 16650 2540 17650 2550
rect 16650 2500 16660 2540
rect 11420 2100 16660 2500
rect 11420 2070 11700 2100
rect 10700 2060 11700 2070
rect 16650 2060 16660 2100
rect 17640 2500 17650 2540
rect 27660 2540 28660 2550
rect 27660 2500 27670 2540
rect 17640 2100 27670 2500
rect 17640 2060 17650 2100
rect 16650 2050 17650 2060
rect 27660 2060 27670 2100
rect 28650 2060 28660 2540
rect 59350 2520 70510 2530
rect 38220 2470 46060 2480
rect 38220 2090 38310 2470
rect 38540 2090 38770 2470
rect 38830 2090 39030 2470
rect 39090 2090 39540 2470
rect 39600 2090 40060 2470
rect 40120 2090 40580 2470
rect 40640 2090 41090 2470
rect 41150 2090 41610 2470
rect 41670 2090 42120 2470
rect 42180 2090 42640 2470
rect 42700 2090 43160 2470
rect 43220 2090 43670 2470
rect 43730 2090 44190 2470
rect 44250 2090 44700 2470
rect 44760 2090 45220 2470
rect 45280 2090 45740 2470
rect 45800 2090 45990 2470
rect 46050 2090 46060 2470
rect 38220 2080 46060 2090
rect 59350 2160 70000 2520
rect 70500 2160 70510 2520
rect 84220 2370 86210 2780
rect 59350 2150 70510 2160
rect 75020 2170 75620 2180
rect 27660 2050 28660 2060
rect 33640 1960 39930 1970
rect 14480 1850 15480 1860
rect 5330 1840 6330 1850
rect 5330 1800 5340 1840
rect 1350 1400 5340 1800
rect 5330 1360 5340 1400
rect 6320 1800 6330 1840
rect 14480 1800 14490 1850
rect 6320 1400 14490 1800
rect 6320 1360 6330 1400
rect 14480 1370 14490 1400
rect 15180 1800 15480 1850
rect 15180 1400 28630 1800
rect 33640 1580 33650 1960
rect 34010 1580 39740 1960
rect 39920 1580 39930 1960
rect 33640 1570 39930 1580
rect 54290 1630 54550 1640
rect 54290 1420 54300 1630
rect 54540 1420 54550 1630
rect 54290 1410 54550 1420
rect 59350 1630 59850 2150
rect 59350 1420 59360 1630
rect 59840 1420 59850 1630
rect 75020 1590 75030 2170
rect 75610 1980 75620 2170
rect 88500 2170 89100 2180
rect 88500 1980 88510 2170
rect 75610 1590 88510 1980
rect 89090 1980 89100 2170
rect 89090 1590 89110 1980
rect 75020 1580 89110 1590
rect 59350 1410 59850 1420
rect 15180 1370 15480 1400
rect 92240 1380 92840 1390
rect 14480 1360 15480 1370
rect 50980 1370 51260 1380
rect 5330 1350 6330 1360
rect 18200 1170 19200 1180
rect 1590 1150 2590 1160
rect 1590 1100 1600 1150
rect 1350 700 1600 1100
rect 1590 670 1600 700
rect 2580 1100 2590 1150
rect 18200 1100 18210 1170
rect 2580 700 18210 1100
rect 2580 670 2590 700
rect 18200 690 18210 700
rect 19190 1100 19200 1170
rect 50980 1110 50990 1370
rect 51250 1350 51260 1370
rect 78800 1370 79400 1380
rect 51250 1130 56760 1350
rect 51250 1110 51260 1130
rect 50980 1100 51260 1110
rect 19190 700 28630 1100
rect 53390 1030 53630 1040
rect 51780 1010 52050 1020
rect 51350 920 51600 930
rect 51350 710 51360 920
rect 51590 710 51600 920
rect 51780 850 51790 1010
rect 52040 850 52050 1010
rect 51780 840 52050 850
rect 53390 840 53400 1030
rect 53620 840 53630 1030
rect 53390 830 53630 840
rect 78800 790 78810 1370
rect 79390 1280 79400 1370
rect 92240 1280 92250 1380
rect 79390 880 92250 1280
rect 79390 790 79400 880
rect 92240 800 92250 880
rect 92830 1280 92840 1380
rect 92830 880 92880 1280
rect 92830 800 92840 880
rect 92240 790 92840 800
rect 78800 780 79400 790
rect 51350 700 51600 710
rect 19190 690 19200 700
rect 18200 680 19200 690
rect 96060 680 96660 690
rect 1590 660 2590 670
rect 82570 670 83170 680
rect 82570 580 82580 670
rect 11340 490 12340 500
rect 7180 390 8780 400
rect 7180 10 7190 390
rect 8770 10 8780 390
rect 7180 0 8780 10
rect 11340 10 11350 490
rect 12330 10 12340 490
rect 11340 0 12340 10
rect 15240 490 16240 500
rect 15240 10 15250 490
rect 16230 10 16240 490
rect 15240 0 16240 10
rect 19460 490 20460 500
rect 19460 10 19470 490
rect 20450 10 20460 490
rect 19460 0 20460 10
rect 22960 490 23960 500
rect 22960 10 22970 490
rect 23950 10 23960 490
rect 22960 0 23960 10
rect 26820 490 27820 500
rect 26820 10 26830 490
rect 27810 10 27820 490
rect 82560 180 82580 580
rect 82570 90 82580 180
rect 83160 580 83170 670
rect 96060 580 96070 680
rect 83160 180 96070 580
rect 83160 90 83170 180
rect 96060 100 96070 180
rect 96650 580 96660 680
rect 96650 180 96670 580
rect 96650 100 96660 180
rect 96060 90 96660 100
rect 82570 80 83170 90
rect 26820 0 27820 10
<< via3 >>
rect 3000 44840 3080 45140
rect 3550 44840 3630 45140
rect 4110 44840 4190 45140
rect 4660 44840 4740 45140
rect 5210 44840 5290 45140
rect 5770 44840 5850 45140
rect 6320 44840 6400 45140
rect 6870 44840 6950 45140
rect 7410 44840 7490 45140
rect 7970 44840 8050 45140
rect 8510 44840 8590 45140
rect 9070 44840 9150 45140
rect 9620 44840 9700 45140
rect 10180 44840 10260 45140
rect 10730 44840 10810 45140
rect 11290 44840 11370 45140
rect 11890 44770 12140 44960
rect 12390 44840 12470 45140
rect 12940 44840 13020 45140
rect 13480 44840 13560 45140
rect 14040 44840 14120 45140
rect 14590 44840 14670 45140
rect 15140 44840 15220 45140
rect 16250 44840 16330 45140
rect 16800 44840 16880 45140
rect 17350 44840 17430 45140
rect 17910 44840 17990 45140
rect 18460 44840 18540 45140
rect 19010 44840 19090 45140
rect 19560 44840 19640 45140
rect 20120 44840 20200 45140
rect 20670 44840 20750 45140
rect 21220 44840 21300 45140
rect 21770 44840 21850 45140
rect 22310 44840 22390 45140
rect 23370 44960 23540 45140
rect 23980 44840 24060 45140
rect 24480 44960 24650 45140
rect 25580 44960 25750 45140
rect 27010 44870 27210 45010
rect 15640 44640 15810 44770
rect 22750 44270 23060 44420
rect 2710 39990 3094 40374
rect 6482 39990 6866 40374
rect 10254 39990 10638 40374
rect 14026 39990 14410 40374
rect 17798 39990 18182 40374
rect 21570 39990 21954 40374
rect 23220 40190 23450 40370
rect 25342 39990 25726 40374
rect 27320 39760 27540 40380
rect 29114 39990 29498 40374
rect 32886 39990 33270 40374
rect 36658 39990 37042 40374
rect 40430 39990 40814 40374
rect 44202 39990 44586 40374
rect 47974 39990 48358 40374
rect 51746 39990 52130 40374
rect 55518 39990 55902 40374
rect 59290 39990 59674 40374
rect 63062 39990 63446 40374
rect 66834 39990 67218 40374
rect 70606 39990 70990 40374
rect 74378 39990 74762 40374
rect 78150 39990 78534 40374
rect 81922 39990 82306 40374
rect 85694 39990 86078 40374
rect 89466 39990 89850 40374
rect 93238 39990 93622 40374
rect 97010 39990 97394 40374
rect 3350 37380 3930 37960
rect 13250 36800 13550 37200
rect 17022 36800 17322 37200
rect 20794 36800 21094 37200
rect 22190 36650 22770 37230
rect 35882 36800 36182 37200
rect 41150 36810 41530 37190
rect 47198 36800 47498 37200
rect 62286 36800 62586 37200
rect 66058 36800 66358 37200
rect 88690 36800 88990 37200
rect 92462 36800 92762 37200
rect 96234 36800 96534 37200
rect 920 36230 1140 36610
rect 4692 36230 4912 36610
rect 8464 36230 8684 36610
rect 12236 36230 12456 36610
rect 16008 36230 16228 36610
rect 19780 36230 20000 36610
rect 23552 36230 23772 36610
rect 27324 36230 27544 36610
rect 31096 36230 31316 36610
rect 34868 36230 35088 36610
rect 38640 36230 38860 36610
rect 42412 36230 42632 36610
rect 46184 36230 46404 36610
rect 49956 36230 50176 36610
rect 53728 36230 53948 36610
rect 57500 36230 57720 36610
rect 61272 36230 61492 36610
rect 65044 36230 65264 36610
rect 68816 36230 69036 36610
rect 72588 36230 72808 36610
rect 76360 36230 76580 36610
rect 80132 36230 80352 36610
rect 83904 36230 84124 36610
rect 87676 36230 87896 36610
rect 91448 36230 91668 36610
rect 95220 36230 95440 36610
rect 2710 35368 3094 35752
rect 6482 35368 6866 35752
rect 10254 35368 10638 35752
rect 14026 35368 14410 35752
rect 17798 35368 18182 35752
rect 21570 35368 21954 35752
rect 23220 35568 23450 35748
rect 25342 35368 25726 35752
rect 27320 35138 27540 35758
rect 29114 35368 29498 35752
rect 32886 35368 33270 35752
rect 36658 35368 37042 35752
rect 40430 35368 40814 35752
rect 44202 35368 44586 35752
rect 47974 35368 48358 35752
rect 51746 35368 52130 35752
rect 55518 35368 55902 35752
rect 59290 35368 59674 35752
rect 63062 35368 63446 35752
rect 66834 35368 67218 35752
rect 70606 35368 70990 35752
rect 74378 35368 74762 35752
rect 78150 35368 78534 35752
rect 81922 35368 82306 35752
rect 85694 35368 86078 35752
rect 89466 35368 89850 35752
rect 93238 35368 93622 35752
rect 97010 35368 97394 35752
rect 7120 32720 7700 33300
rect 13250 32178 13550 32578
rect 17022 32178 17322 32578
rect 20794 32178 21094 32578
rect 25980 32030 26560 32610
rect 35882 32178 36182 32578
rect 47198 32178 47498 32578
rect 48700 32190 49070 32570
rect 62286 32178 62586 32578
rect 66058 32178 66358 32578
rect 88690 32178 88990 32578
rect 92462 32178 92762 32578
rect 96234 32178 96534 32578
rect 2710 30746 3094 31130
rect 6482 30746 6866 31130
rect 10254 30746 10638 31130
rect 14026 30746 14410 31130
rect 17798 30746 18182 31130
rect 21570 30746 21954 31130
rect 23220 30946 23450 31126
rect 25342 30746 25726 31130
rect 27320 30516 27540 31136
rect 29114 30746 29498 31130
rect 32886 30746 33270 31130
rect 36658 30746 37042 31130
rect 40430 30746 40814 31130
rect 44202 30746 44586 31130
rect 47974 30746 48358 31130
rect 51746 30746 52130 31130
rect 55518 30746 55902 31130
rect 59290 30746 59674 31130
rect 63062 30746 63446 31130
rect 66834 30746 67218 31130
rect 70606 30746 70990 31130
rect 74378 30746 74762 31130
rect 78150 30746 78534 31130
rect 81922 30746 82306 31130
rect 85694 30746 86078 31130
rect 89466 30746 89850 31130
rect 93238 30746 93622 31130
rect 97010 30746 97394 31130
rect 10900 28100 11480 28680
rect 13250 27556 13550 27956
rect 17022 27556 17322 27956
rect 20794 27556 21094 27956
rect 29730 27440 30310 28020
rect 35882 27556 36182 27956
rect 47198 27556 47498 27956
rect 56240 27570 56620 27940
rect 62286 27556 62586 27956
rect 66058 27556 66358 27956
rect 88690 27556 88990 27956
rect 92462 27556 92762 27956
rect 96234 27556 96534 27956
rect 2710 26124 3094 26508
rect 6482 26124 6866 26508
rect 10254 26124 10638 26508
rect 14026 26124 14410 26508
rect 17798 26124 18182 26508
rect 21570 26124 21954 26508
rect 23220 26324 23450 26504
rect 25342 26124 25726 26508
rect 27320 25894 27540 26514
rect 29114 26124 29498 26508
rect 32886 26124 33270 26508
rect 36658 26124 37042 26508
rect 40430 26124 40814 26508
rect 44802 26124 45186 26508
rect 47974 26124 48358 26508
rect 52346 26124 52730 26508
rect 55518 26124 55902 26508
rect 59290 26124 59674 26508
rect 63062 26124 63446 26508
rect 66834 26124 67218 26508
rect 71206 26124 71590 26508
rect 74378 26124 74762 26508
rect 78150 26124 78534 26508
rect 81922 26124 82306 26508
rect 85694 26124 86078 26508
rect 89466 26124 89850 26508
rect 93238 26124 93622 26508
rect 97010 26124 97394 26508
rect 14670 23480 15250 24060
rect 90140 23470 90650 24150
rect 13250 22934 13550 23334
rect 17022 22934 17322 23334
rect 20794 22934 21094 23334
rect 35882 22934 36182 23334
rect 47198 22934 47498 23334
rect 62286 22934 62586 23334
rect 66058 22934 66358 23334
rect 41150 22350 41530 22730
rect 43426 22340 43726 22740
rect 50970 22340 51270 22740
rect 69830 22340 70130 22740
rect 75130 22390 75520 23370
rect 88690 22934 88990 23334
rect 92462 22934 92762 23334
rect 96234 22934 96534 23334
rect 2710 21502 3094 21886
rect 6482 21502 6866 21886
rect 10254 21502 10638 21886
rect 14026 21502 14410 21886
rect 17798 21502 18182 21886
rect 21570 21502 21954 21886
rect 23220 21702 23450 21882
rect 25342 21502 25726 21886
rect 27320 21272 27540 21892
rect 29114 21502 29498 21886
rect 32886 21502 33270 21886
rect 36658 21502 37042 21886
rect 40430 21502 40814 21886
rect 44802 21502 45186 21886
rect 47974 21502 48358 21886
rect 52346 21502 52730 21886
rect 55518 21502 55902 21886
rect 59290 21502 59674 21886
rect 63062 21502 63446 21886
rect 66834 21502 67218 21886
rect 71206 21502 71590 21886
rect 74378 21502 74762 21886
rect 78150 21502 78534 21886
rect 81922 21502 82306 21886
rect 85694 21502 86078 21886
rect 89466 21502 89850 21886
rect 93238 21502 93622 21886
rect 97010 21502 97394 21886
rect 18430 18860 19010 19440
rect 93910 18840 94420 19520
rect 13250 18312 13550 18712
rect 17022 18312 17322 18712
rect 20794 18312 21094 18712
rect 35882 18312 36182 18712
rect 47198 18312 47498 18712
rect 62286 18312 62586 18712
rect 66058 18312 66358 18712
rect 43426 17718 43726 18118
rect 48700 17730 49070 18110
rect 50970 17718 51270 18118
rect 69830 17718 70130 18118
rect 78910 17760 79290 18740
rect 88690 18312 88990 18712
rect 92462 18312 92762 18712
rect 96234 18312 96534 18712
rect 2710 16880 3094 17264
rect 6482 16880 6866 17264
rect 10254 16880 10638 17264
rect 14026 16880 14410 17264
rect 17798 16880 18182 17264
rect 21570 16880 21954 17264
rect 23220 17080 23450 17260
rect 25342 16880 25726 17264
rect 27320 16650 27540 17270
rect 29114 16880 29498 17264
rect 32886 16880 33270 17264
rect 36658 16880 37042 17264
rect 40430 16880 40814 17264
rect 44802 16880 45186 17264
rect 47974 16880 48358 17264
rect 52346 16880 52730 17264
rect 55518 16880 55902 17264
rect 59290 16880 59674 17264
rect 63062 16880 63446 17264
rect 66834 16880 67218 17264
rect 71206 16880 71590 17264
rect 74378 16880 74762 17264
rect 78150 16880 78534 17264
rect 81922 16880 82306 17264
rect 85694 16880 86078 17264
rect 89466 16880 89850 17264
rect 93238 16880 93622 17264
rect 97010 16880 97394 17264
rect 13250 13690 13550 14090
rect 17022 13690 17322 14090
rect 20794 13690 21094 14090
rect 35882 13690 36182 14090
rect 47198 13690 47498 14090
rect 62286 13690 62586 14090
rect 66058 13690 66358 14090
rect 43426 13096 43726 13496
rect 50970 13096 51270 13496
rect 56240 13110 56610 13480
rect 69830 13096 70130 13496
rect 82680 13110 83060 14090
rect 88690 13690 88990 14090
rect 92462 13690 92762 14090
rect 96234 13690 96534 14090
rect 97770 13700 98150 14680
rect 10250 12260 10640 12650
rect 14020 12260 14410 12650
rect 25270 12260 25850 12840
rect 29090 12260 29670 12840
rect 70610 12770 70980 12960
rect 71210 12500 71580 12690
rect 85700 12270 86070 12640
rect 89470 12270 89840 12640
rect 66840 11050 67210 11430
rect 2710 10560 3090 10940
rect 8130 10550 8370 10940
rect 11900 10550 12140 10940
rect 32880 10550 33270 10940
rect 33650 10430 34020 10930
rect 36650 10550 37040 10940
rect 37420 10430 37790 10930
rect 59290 10560 59670 10940
rect 63060 10560 63440 10940
rect 78150 10560 78530 10940
rect 83580 10570 83800 10930
rect 87350 10560 87570 10940
rect 97010 10560 97390 10940
rect 22330 9340 22710 10030
rect 26090 9370 26470 10060
rect 70610 9940 70980 10130
rect 74380 10020 74750 10410
rect 71210 9670 71580 9860
rect 86530 8960 86880 9340
rect 8460 7710 8680 8180
rect 12230 7720 12450 8180
rect 29720 8190 30300 8780
rect 63060 8160 63440 8480
rect 81920 8350 82300 8590
rect 47980 7670 48350 8050
rect 44800 7030 45180 7410
rect 52340 7230 52720 7610
rect 90220 7300 90600 8020
rect 94000 7300 94380 8020
rect 97770 7300 98150 8020
rect 10250 5590 10640 6350
rect 46180 6410 46430 6790
rect 14020 5590 14410 6350
rect 32880 5930 33270 6320
rect 36650 5930 37040 6320
rect 6480 5130 6860 5310
rect 2710 4810 3090 4990
rect 38630 5420 38860 6040
rect 40430 5760 40810 5940
rect 44200 5810 44580 6190
rect 51740 5810 52120 6190
rect 59290 5930 59670 6320
rect 63060 5930 63440 6320
rect 85690 6190 85820 6580
rect 85820 6190 85880 6580
rect 85880 6190 86070 6580
rect 40430 5560 40810 5760
rect 50660 5390 50880 5680
rect 55520 5390 55900 5740
rect 17790 5120 18180 5320
rect 21570 4800 21950 5000
rect 37420 4870 37790 5250
rect 78150 5210 78530 5550
rect 36650 4340 37040 4720
rect 3150 3410 3860 3890
rect 24060 3470 25040 3950
rect 33650 3850 34020 4230
rect 50660 3830 50880 4210
rect 51010 4070 51230 4460
rect 86530 4590 86880 4960
rect 38310 3310 38540 3690
rect 46180 3250 46610 3630
rect 6910 2770 7620 3250
rect 20440 2760 21420 3240
rect 28870 2760 29850 3240
rect 32880 2610 33270 2990
rect 59300 2860 59660 3500
rect 65040 3220 65480 3800
rect 97010 3530 97390 3930
rect 89470 2870 89840 3260
rect 93240 2870 93620 3260
rect 10710 2070 11420 2550
rect 16660 2060 17640 2540
rect 27670 2060 28650 2540
rect 38310 2090 38540 2470
rect 5340 1360 6320 1840
rect 14490 1370 15180 1850
rect 54300 1420 54540 1630
rect 59360 1420 59840 1630
rect 75030 1590 75610 2170
rect 88510 1590 89090 2170
rect 1600 670 2580 1150
rect 18210 690 19190 1170
rect 50990 1110 51250 1370
rect 51360 710 51590 920
rect 51790 850 52040 1010
rect 53400 840 53620 1030
rect 78810 790 79390 1370
rect 92250 800 92830 1380
rect 7190 10 8770 390
rect 11350 10 12330 490
rect 15250 10 16230 490
rect 19470 10 20450 490
rect 22970 10 23950 490
rect 26830 10 27810 490
rect 82580 90 83160 670
rect 96070 100 96650 680
<< metal4 >>
rect 3006 45150 3066 45152
rect 3558 45150 3618 45152
rect 4110 45150 4170 45152
rect 4662 45150 4722 45152
rect 5214 45150 5274 45152
rect 5766 45150 5826 45152
rect 6318 45150 6378 45152
rect 6870 45150 6930 45152
rect 7422 45150 7482 45152
rect 7974 45150 8034 45152
rect 8526 45150 8586 45152
rect 9078 45150 9138 45152
rect 9630 45150 9690 45152
rect 10182 45150 10242 45152
rect 10734 45150 10794 45152
rect 11286 45150 11346 45152
rect 11838 45150 11898 45152
rect 12390 45150 12450 45152
rect 12942 45150 13002 45152
rect 13494 45150 13554 45152
rect 14046 45150 14106 45152
rect 14598 45150 14658 45152
rect 15150 45150 15210 45152
rect 15702 45150 15762 45152
rect 16254 45150 16314 45152
rect 16806 45150 16866 45152
rect 17358 45150 17418 45152
rect 17910 45150 17970 45152
rect 18462 45150 18522 45152
rect 19014 45150 19074 45152
rect 19566 45150 19626 45152
rect 20118 45150 20178 45152
rect 20670 45150 20730 45152
rect 21222 45150 21282 45152
rect 21774 45150 21834 45152
rect 22326 45150 22386 45152
rect 22878 45150 22938 45152
rect 23430 45150 23490 45152
rect 23982 45150 24042 45152
rect 24534 45150 24594 45152
rect 2990 45140 3090 45150
rect 2990 44840 3000 45140
rect 3080 44840 3090 45140
rect 2990 44830 3090 44840
rect 3540 45140 3640 45150
rect 3540 44840 3550 45140
rect 3630 44840 3640 45140
rect 3540 44830 3640 44840
rect 4100 45140 4200 45150
rect 4100 44840 4110 45140
rect 4190 44840 4200 45140
rect 4100 44830 4200 44840
rect 4650 45140 4750 45150
rect 4650 44840 4660 45140
rect 4740 44840 4750 45140
rect 4650 44830 4750 44840
rect 5200 45140 5300 45150
rect 5200 44840 5210 45140
rect 5290 44840 5300 45140
rect 5200 44830 5300 44840
rect 5760 45140 5860 45150
rect 5760 44840 5770 45140
rect 5850 44840 5860 45140
rect 5760 44830 5860 44840
rect 6310 45140 6410 45150
rect 6310 44840 6320 45140
rect 6400 44840 6410 45140
rect 6310 44830 6410 44840
rect 6860 45140 6960 45150
rect 6860 44840 6870 45140
rect 6950 44840 6960 45140
rect 6860 44830 6960 44840
rect 7400 45140 7500 45150
rect 7400 44840 7410 45140
rect 7490 44840 7500 45140
rect 7400 44830 7500 44840
rect 7960 45140 8060 45150
rect 7960 44840 7970 45140
rect 8050 44840 8060 45140
rect 7960 44830 8060 44840
rect 8500 45140 8600 45150
rect 8500 44840 8510 45140
rect 8590 44840 8600 45140
rect 8500 44830 8600 44840
rect 9060 45140 9160 45150
rect 9060 44840 9070 45140
rect 9150 44840 9160 45140
rect 9060 44830 9160 44840
rect 9610 45140 9710 45150
rect 9610 44840 9620 45140
rect 9700 44840 9710 45140
rect 9610 44830 9710 44840
rect 10170 45140 10270 45150
rect 10170 44840 10180 45140
rect 10260 44840 10270 45140
rect 10170 44830 10270 44840
rect 10720 45140 10820 45150
rect 10720 44840 10730 45140
rect 10810 44840 10820 45140
rect 10720 44830 10820 44840
rect 11280 45140 11380 45150
rect 11280 44840 11290 45140
rect 11370 44840 11380 45140
rect 11280 44830 11380 44840
rect 11820 44970 11920 45150
rect 12380 45140 12480 45150
rect 11820 44960 12150 44970
rect 11820 44830 11890 44960
rect 11880 44770 11890 44830
rect 12140 44770 12150 44960
rect 12380 44840 12390 45140
rect 12470 44840 12480 45140
rect 12380 44830 12480 44840
rect 12930 45140 13030 45150
rect 12930 44840 12940 45140
rect 13020 44840 13030 45140
rect 12930 44830 13030 44840
rect 13470 45140 13570 45150
rect 13470 44840 13480 45140
rect 13560 44840 13570 45140
rect 13470 44830 13570 44840
rect 14030 45140 14130 45150
rect 14030 44840 14040 45140
rect 14120 44840 14130 45140
rect 14030 44830 14130 44840
rect 14580 45140 14680 45150
rect 14580 44840 14590 45140
rect 14670 44840 14680 45140
rect 14580 44830 14680 44840
rect 15130 45140 15230 45150
rect 15130 44840 15140 45140
rect 15220 44840 15230 45140
rect 15130 44830 15230 44840
rect 11880 44760 12150 44770
rect 15630 44770 15820 45150
rect 16240 45140 16340 45150
rect 16240 44840 16250 45140
rect 16330 44840 16340 45140
rect 16240 44830 16340 44840
rect 16790 45140 16890 45150
rect 16790 44840 16800 45140
rect 16880 44840 16890 45140
rect 16790 44830 16890 44840
rect 17340 45140 17440 45150
rect 17340 44840 17350 45140
rect 17430 44840 17440 45140
rect 17340 44830 17440 44840
rect 17900 45140 18000 45150
rect 17900 44840 17910 45140
rect 17990 44840 18000 45140
rect 17900 44830 18000 44840
rect 18450 45140 18550 45150
rect 18450 44840 18460 45140
rect 18540 44840 18550 45140
rect 18450 44830 18550 44840
rect 19000 45140 19100 45150
rect 19000 44840 19010 45140
rect 19090 44840 19100 45140
rect 19000 44830 19100 44840
rect 19550 45140 19650 45150
rect 19550 44840 19560 45140
rect 19640 44840 19650 45140
rect 19550 44830 19650 44840
rect 20110 45140 20210 45150
rect 20110 44840 20120 45140
rect 20200 44840 20210 45140
rect 20110 44830 20210 44840
rect 20660 45140 20760 45150
rect 20660 44840 20670 45140
rect 20750 44840 20760 45140
rect 20660 44830 20760 44840
rect 21210 45140 21310 45150
rect 21210 44840 21220 45140
rect 21300 44840 21310 45140
rect 21210 44830 21310 44840
rect 21760 45140 21860 45150
rect 21760 44840 21770 45140
rect 21850 44840 21860 45140
rect 21760 44830 21860 44840
rect 22300 45140 22400 45150
rect 22300 44840 22310 45140
rect 22390 44840 22400 45140
rect 22300 44830 22400 44840
rect 300 43980 480 44160
rect 620 43980 800 44160
rect 940 43980 1120 44160
rect 11910 44080 12120 44760
rect 15630 44640 15640 44770
rect 15810 44640 15820 44770
rect 15630 44630 15820 44640
rect 22810 44430 23000 45150
rect 23360 45140 23550 45150
rect 23360 44960 23370 45140
rect 23540 44960 23550 45140
rect 23360 44950 23550 44960
rect 23970 45140 24070 45150
rect 23970 44840 23980 45140
rect 24060 44840 24070 45140
rect 24470 45140 24660 45150
rect 24470 44960 24480 45140
rect 24650 44960 24660 45140
rect 24470 44950 24660 44960
rect 25086 44952 25146 45152
rect 25638 45150 25698 45152
rect 25570 45140 25760 45150
rect 25570 44960 25580 45140
rect 25750 44960 25760 45140
rect 25570 44950 25760 44960
rect 26190 44952 26250 45152
rect 27000 45010 27220 45020
rect 23970 44830 24070 44840
rect 27000 44870 27010 45010
rect 27210 44870 27220 45010
rect 22740 44420 23070 44430
rect 22740 44270 22750 44420
rect 23060 44270 23070 44420
rect 22740 44260 23070 44270
rect 27000 44050 27220 44870
rect 2700 40374 3100 40600
rect 2700 39990 2710 40374
rect 3094 39990 3100 40374
rect 2700 35752 3100 39990
rect 6472 40374 6872 40600
rect 6472 39990 6482 40374
rect 6866 39990 6872 40374
rect 3340 37960 3940 37970
rect 3340 37380 3350 37960
rect 3930 37380 3940 37960
rect 3340 37370 3940 37380
rect 2700 35368 2710 35752
rect 3094 35368 3100 35752
rect 2700 31130 3100 35368
rect 2700 30746 2710 31130
rect 3094 30746 3100 31130
rect 2700 26508 3100 30746
rect 2700 26124 2710 26508
rect 3094 26124 3100 26508
rect 2700 21886 3100 26124
rect 2700 21502 2710 21886
rect 3094 21502 3100 21886
rect 2700 17264 3100 21502
rect 2700 16880 2710 17264
rect 3094 16880 3100 17264
rect 2700 10940 3100 16880
rect 2700 10560 2710 10940
rect 3090 10560 3100 10940
rect 1890 1160 2290 6920
rect 2700 4990 3100 10560
rect 2700 4810 2710 4990
rect 3090 4810 3100 4990
rect 2700 4790 3100 4810
rect 3460 3900 3860 37370
rect 6472 35752 6872 39990
rect 10244 40374 10644 40600
rect 10244 39990 10254 40374
rect 10638 39990 10644 40374
rect 6472 35368 6482 35752
rect 6866 35368 6872 35752
rect 6472 31130 6872 35368
rect 10244 35752 10644 39990
rect 14016 40374 14416 40600
rect 14016 39990 14026 40374
rect 14410 39990 14416 40374
rect 13300 37210 13500 39090
rect 13240 37200 13560 37210
rect 13240 36800 13250 37200
rect 13550 36800 13560 37200
rect 13240 36790 13560 36800
rect 10244 35368 10254 35752
rect 10638 35368 10644 35752
rect 7110 33300 7710 33310
rect 7110 32720 7120 33300
rect 7700 32720 7710 33300
rect 7110 32710 7710 32720
rect 6472 30746 6482 31130
rect 6866 30746 6872 31130
rect 6472 26508 6872 30746
rect 6472 26124 6482 26508
rect 6866 26124 6872 26508
rect 6472 21886 6872 26124
rect 6472 21502 6482 21886
rect 6866 21502 6872 21886
rect 6472 17264 6872 21502
rect 6472 16880 6482 17264
rect 6866 16880 6872 17264
rect 3140 3890 3880 3900
rect 3140 3410 3150 3890
rect 3860 3410 3880 3890
rect 3140 3400 3880 3410
rect 5660 1850 6060 6930
rect 6472 5310 6872 16880
rect 6472 5130 6480 5310
rect 6860 5130 6872 5310
rect 6472 5120 6872 5130
rect 7220 3260 7620 32710
rect 10244 31130 10644 35368
rect 14016 35752 14416 39990
rect 17788 40374 18188 40600
rect 17788 39990 17798 40374
rect 18182 39990 18188 40374
rect 17072 37210 17272 39090
rect 17012 37200 17332 37210
rect 17012 36800 17022 37200
rect 17322 36800 17332 37200
rect 17012 36790 17332 36800
rect 14016 35368 14026 35752
rect 14410 35368 14416 35752
rect 13300 32588 13500 34468
rect 13240 32578 13560 32588
rect 13240 32178 13250 32578
rect 13550 32178 13560 32578
rect 13240 32168 13560 32178
rect 10244 30746 10254 31130
rect 10638 30746 10644 31130
rect 10244 26508 10644 30746
rect 14016 31130 14416 35368
rect 17788 35752 18188 39990
rect 21560 40374 21960 40600
rect 21560 39990 21570 40374
rect 21954 39990 21960 40374
rect 25332 40374 25732 40600
rect 20844 37210 21044 39090
rect 20784 37200 21104 37210
rect 20784 36800 20794 37200
rect 21094 36800 21104 37200
rect 20784 36790 21104 36800
rect 17788 35368 17798 35752
rect 18182 35368 18188 35752
rect 17072 32588 17272 34468
rect 17012 32578 17332 32588
rect 17012 32178 17022 32578
rect 17322 32178 17332 32578
rect 17012 32168 17332 32178
rect 14016 30746 14026 31130
rect 14410 30746 14416 31130
rect 10890 28680 11490 28690
rect 10890 28100 10900 28680
rect 11480 28100 11490 28680
rect 10890 28090 11490 28100
rect 10244 26124 10254 26508
rect 10638 26124 10644 26508
rect 10244 21886 10644 26124
rect 10244 21502 10254 21886
rect 10638 21502 10644 21886
rect 10244 17264 10644 21502
rect 10244 16880 10254 17264
rect 10638 16880 10644 17264
rect 10244 12650 10644 16880
rect 10244 12260 10250 12650
rect 10640 12260 10644 12650
rect 8120 10940 8380 10960
rect 8120 10550 8130 10940
rect 8370 10550 8380 10940
rect 8120 10540 8380 10550
rect 10244 6350 10644 12260
rect 10244 5590 10250 6350
rect 10640 5590 10644 6350
rect 10244 5580 10644 5590
rect 6900 3250 7640 3260
rect 6900 2770 6910 3250
rect 7620 2770 7640 3250
rect 6900 2760 7640 2770
rect 11010 2560 11410 28090
rect 13300 27966 13500 29846
rect 13240 27956 13560 27966
rect 13240 27556 13250 27956
rect 13550 27556 13560 27956
rect 13240 27546 13560 27556
rect 14016 26508 14416 30746
rect 17788 31130 18188 35368
rect 21560 35752 21960 39990
rect 25332 39990 25342 40374
rect 25726 39990 25732 40374
rect 22180 37230 22780 37240
rect 22180 36650 22190 37230
rect 22770 36650 22780 37230
rect 22180 36640 22780 36650
rect 21560 35368 21570 35752
rect 21954 35368 21960 35752
rect 20844 32588 21044 34468
rect 20784 32578 21104 32588
rect 20784 32178 20794 32578
rect 21094 32178 21104 32578
rect 20784 32168 21104 32178
rect 17788 30746 17798 31130
rect 18182 30746 18188 31130
rect 17072 27966 17272 29846
rect 17012 27956 17332 27966
rect 17012 27556 17022 27956
rect 17322 27556 17332 27956
rect 17012 27546 17332 27556
rect 14016 26124 14026 26508
rect 14410 26124 14416 26508
rect 13300 23344 13500 25224
rect 13240 23334 13560 23344
rect 13240 22934 13250 23334
rect 13550 22934 13560 23334
rect 13240 22924 13560 22934
rect 14016 21886 14416 26124
rect 17788 26508 18188 30746
rect 21560 31130 21960 35368
rect 21560 30746 21570 31130
rect 21954 30746 21960 31130
rect 20844 27966 21044 29846
rect 20784 27956 21104 27966
rect 20784 27556 20794 27956
rect 21094 27556 21104 27956
rect 20784 27546 21104 27556
rect 17788 26124 17798 26508
rect 18182 26124 18188 26508
rect 14660 24060 15260 24070
rect 14660 23480 14670 24060
rect 15250 23480 15260 24060
rect 14660 23470 15260 23480
rect 14016 21502 14026 21886
rect 14410 21502 14416 21886
rect 13300 18722 13500 20602
rect 13240 18712 13560 18722
rect 13240 18312 13250 18712
rect 13550 18312 13560 18712
rect 13240 18302 13560 18312
rect 14016 17264 14416 21502
rect 14016 16880 14026 17264
rect 14410 16880 14416 17264
rect 13300 14100 13500 15980
rect 13240 14090 13560 14100
rect 13240 13690 13250 14090
rect 13550 13690 13560 14090
rect 13240 13680 13560 13690
rect 14016 12650 14416 16880
rect 14016 12260 14020 12650
rect 14410 12260 14416 12650
rect 11890 10940 12150 10960
rect 11890 10550 11900 10940
rect 12140 10550 12150 10940
rect 11890 10540 12150 10550
rect 14016 6350 14416 12260
rect 14016 5590 14020 6350
rect 14410 5590 14416 6350
rect 14016 5560 14416 5590
rect 10700 2550 11440 2560
rect 10700 2070 10710 2550
rect 11420 2070 11440 2550
rect 10700 2060 11440 2070
rect 14780 1860 15180 23470
rect 17072 23344 17272 25224
rect 17012 23334 17332 23344
rect 17012 22934 17022 23334
rect 17322 22934 17332 23334
rect 17012 22924 17332 22934
rect 17788 21886 18188 26124
rect 21560 26508 21960 30746
rect 21560 26124 21570 26508
rect 21954 26124 21960 26508
rect 20844 23344 21044 25224
rect 20784 23334 21104 23344
rect 20784 22934 20794 23334
rect 21094 22934 21104 23334
rect 20784 22924 21104 22934
rect 17788 21502 17798 21886
rect 18182 21502 18188 21886
rect 17072 18722 17272 20602
rect 17012 18712 17332 18722
rect 17012 18312 17022 18712
rect 17322 18312 17332 18712
rect 17012 18302 17332 18312
rect 17788 17264 18188 21502
rect 21560 21886 21960 26124
rect 21560 21502 21570 21886
rect 21954 21502 21960 21886
rect 18420 19440 19020 19450
rect 18420 18860 18430 19440
rect 19010 18860 19020 19440
rect 18420 18850 19020 18860
rect 17788 16880 17798 17264
rect 18182 16880 18188 17264
rect 17072 14100 17272 15980
rect 17012 14090 17332 14100
rect 17012 13690 17022 14090
rect 17322 13690 17332 14090
rect 17012 13680 17332 13690
rect 16970 2550 17370 6840
rect 17788 5320 18188 16880
rect 18550 5710 18950 18850
rect 20844 18722 21044 20602
rect 20784 18712 21104 18722
rect 20784 18312 20794 18712
rect 21094 18312 21104 18712
rect 20784 18302 21104 18312
rect 21560 17264 21960 21502
rect 21560 16880 21570 17264
rect 21954 16880 21960 17264
rect 20844 14100 21044 15980
rect 20784 14090 21104 14100
rect 20784 13690 20794 14090
rect 21094 13690 21104 14090
rect 20784 13680 21104 13690
rect 17788 5120 17790 5320
rect 18180 5120 18188 5320
rect 17788 5090 18188 5120
rect 18510 5110 18980 5710
rect 16650 2540 17650 2550
rect 16650 2060 16660 2540
rect 17640 2060 17650 2540
rect 16650 2050 17650 2060
rect 14480 1850 15190 1860
rect 5330 1840 6330 1850
rect 5330 1360 5340 1840
rect 6320 1360 6330 1840
rect 14480 1370 14490 1850
rect 15180 1370 15190 1850
rect 14480 1360 15190 1370
rect 5330 1350 6330 1360
rect 18550 1180 18950 5110
rect 20740 3250 21140 6820
rect 21560 5000 21960 16880
rect 22320 10030 22720 36640
rect 25332 35752 25732 39990
rect 29104 40374 29504 40600
rect 29104 39990 29114 40374
rect 29498 39990 29504 40374
rect 25332 35368 25342 35752
rect 25726 35368 25732 35752
rect 25332 31130 25732 35368
rect 29104 35752 29504 39990
rect 32876 40374 33276 40600
rect 32876 39990 32886 40374
rect 33270 39990 33276 40374
rect 29104 35368 29114 35752
rect 29498 35368 29504 35752
rect 26080 32620 26480 32700
rect 25970 32610 26570 32620
rect 25970 32030 25980 32610
rect 26560 32030 26570 32610
rect 25970 32020 26570 32030
rect 25332 30746 25342 31130
rect 25726 30746 25732 31130
rect 25332 26508 25732 30746
rect 25332 26124 25342 26508
rect 25726 26124 25732 26508
rect 25332 21886 25732 26124
rect 25332 21502 25342 21886
rect 25726 21502 25732 21886
rect 25332 17264 25732 21502
rect 25332 16880 25342 17264
rect 25726 16880 25732 17264
rect 25332 16000 25732 16880
rect 25260 12840 25860 12850
rect 25260 12260 25270 12840
rect 25850 12260 25860 12840
rect 25260 12250 25860 12260
rect 22320 9340 22330 10030
rect 22710 9340 22720 10030
rect 22320 9330 22720 9340
rect 25350 6830 25750 12250
rect 26080 10060 26480 32020
rect 29104 31130 29504 35368
rect 29104 30746 29114 31130
rect 29498 30746 29504 31130
rect 29104 26508 29504 30746
rect 32876 35752 33276 39990
rect 36648 40374 37048 40600
rect 36648 39990 36658 40374
rect 37042 39990 37048 40374
rect 35932 37210 36132 39090
rect 35870 37200 36190 37210
rect 35870 36800 35882 37200
rect 36182 36800 36190 37200
rect 35870 36790 36190 36800
rect 32876 35368 32886 35752
rect 33270 35368 33276 35752
rect 32876 31130 33276 35368
rect 36648 35752 37048 39990
rect 40420 40374 40820 40600
rect 40420 39990 40430 40374
rect 40814 39990 40820 40374
rect 36648 35368 36658 35752
rect 37042 35368 37048 35752
rect 35932 32588 36132 34468
rect 35870 32578 36190 32588
rect 35870 32178 35882 32578
rect 36182 32178 36190 32578
rect 35870 32168 36190 32178
rect 32876 30746 32886 31130
rect 33270 30746 33276 31130
rect 29860 28030 30260 28060
rect 29720 28020 30320 28030
rect 29720 27440 29730 28020
rect 30310 27440 30320 28020
rect 29720 27430 30320 27440
rect 29104 26124 29114 26508
rect 29498 26124 29504 26508
rect 29104 21886 29504 26124
rect 29104 21502 29114 21886
rect 29498 21502 29504 21886
rect 29104 17264 29504 21502
rect 29104 16880 29114 17264
rect 29498 16880 29504 17264
rect 29104 16000 29504 16880
rect 29080 12840 29680 12850
rect 29080 12260 29090 12840
rect 29670 12260 29680 12840
rect 29080 12250 29680 12260
rect 26080 9370 26090 10060
rect 26470 9370 26480 10060
rect 26080 9360 26480 9370
rect 21560 4800 21570 5000
rect 21950 4800 21960 5000
rect 21560 4730 21960 4800
rect 24510 6250 25750 6830
rect 24510 3960 24910 6250
rect 24050 3950 25050 3960
rect 24050 3470 24060 3950
rect 25040 3470 25050 3950
rect 24050 3460 25050 3470
rect 29110 3250 29510 12250
rect 29860 8790 30260 27430
rect 32876 26508 33276 30746
rect 36648 31130 37048 35368
rect 36648 30746 36658 31130
rect 37042 30746 37048 31130
rect 35932 27966 36132 29846
rect 35870 27956 36190 27966
rect 35870 27556 35882 27956
rect 36182 27556 36190 27956
rect 35870 27546 36190 27556
rect 32876 26124 32886 26508
rect 33270 26124 33276 26508
rect 32876 21886 33276 26124
rect 36648 26508 37048 30746
rect 36648 26124 36658 26508
rect 37042 26124 37048 26508
rect 35932 23344 36132 25224
rect 35870 23334 36190 23344
rect 35870 22934 35882 23334
rect 36182 22934 36190 23334
rect 35870 22924 36190 22934
rect 32876 21502 32886 21886
rect 33270 21502 33276 21886
rect 32876 17264 33276 21502
rect 36648 21886 37048 26124
rect 36648 21502 36658 21886
rect 37042 21502 37048 21886
rect 35932 18722 36132 20602
rect 35870 18712 36190 18722
rect 35870 18312 35882 18712
rect 36182 18312 36190 18712
rect 35870 18302 36190 18312
rect 32876 16880 32886 17264
rect 33270 16880 33276 17264
rect 32876 16000 33276 16880
rect 36648 17264 37048 21502
rect 36648 16880 36658 17264
rect 37042 16880 37048 17264
rect 36648 16000 37048 16880
rect 40420 35752 40820 39990
rect 44192 40374 44592 40600
rect 44192 39990 44202 40374
rect 44586 39990 44592 40374
rect 40420 35368 40430 35752
rect 40814 35368 40820 35752
rect 40420 31130 40820 35368
rect 40420 30746 40430 31130
rect 40814 30746 40820 31130
rect 40420 26508 40820 30746
rect 40420 26124 40430 26508
rect 40814 26124 40820 26508
rect 40420 21886 40820 26124
rect 41140 37190 41540 37810
rect 41140 36810 41150 37190
rect 41530 36810 41540 37190
rect 41140 22730 41540 36810
rect 44192 35752 44592 39990
rect 44192 35368 44202 35752
rect 44586 35368 44592 35752
rect 44192 31130 44592 35368
rect 44192 30746 44202 31130
rect 44586 30746 44592 31130
rect 43476 22750 43676 25224
rect 41140 22350 41150 22730
rect 41530 22350 41540 22730
rect 41140 22340 41540 22350
rect 43414 22740 43734 22750
rect 43414 22340 43426 22740
rect 43726 22340 43734 22740
rect 43414 22330 43734 22340
rect 40420 21502 40430 21886
rect 40814 21502 40820 21886
rect 40420 17264 40820 21502
rect 43476 18128 43676 20602
rect 43414 18118 43734 18128
rect 43414 17718 43426 18118
rect 43726 17718 43734 18118
rect 43414 17708 43734 17718
rect 40420 16880 40430 17264
rect 40814 16880 40820 17264
rect 32870 10940 33280 16000
rect 35932 14100 36132 15980
rect 35870 14090 36190 14100
rect 35870 13690 35882 14090
rect 36182 13690 36190 14090
rect 35870 13680 36190 13690
rect 36640 10940 37050 16000
rect 32870 10550 32880 10940
rect 33270 10550 33280 10940
rect 29710 8780 30310 8790
rect 29710 8190 29720 8780
rect 30300 8190 30310 8780
rect 29710 8180 30310 8190
rect 32870 6320 33280 10550
rect 32870 5930 32880 6320
rect 33270 5930 33280 6320
rect 20430 3240 21430 3250
rect 20430 2760 20440 3240
rect 21420 2760 21430 3240
rect 20430 2750 21430 2760
rect 28860 3240 29860 3250
rect 28860 2760 28870 3240
rect 29850 2760 29860 3240
rect 28860 2750 29860 2760
rect 32870 2990 33280 5930
rect 33640 10930 34030 10940
rect 33640 10430 33650 10930
rect 34020 10430 34030 10930
rect 33640 4230 34030 10430
rect 33640 3850 33650 4230
rect 34020 3850 34030 4230
rect 33640 3840 34030 3850
rect 36640 10550 36650 10940
rect 37040 10550 37050 10940
rect 36640 6320 37050 10550
rect 36640 5930 36650 6320
rect 37040 5930 37050 6320
rect 36640 4720 37050 5930
rect 37410 10930 37800 10940
rect 37410 10430 37420 10930
rect 37790 10430 37800 10930
rect 37410 5250 37800 10430
rect 38620 6040 38870 6050
rect 38620 5420 38630 6040
rect 38860 5420 38870 6040
rect 40420 5940 40820 16880
rect 43476 13506 43676 15980
rect 43414 13496 43734 13506
rect 43414 13096 43426 13496
rect 43726 13096 43734 13496
rect 43414 13086 43734 13096
rect 44192 6200 44592 30746
rect 44792 26508 45192 40600
rect 47964 40374 48364 40600
rect 47964 39990 47974 40374
rect 48358 39990 48364 40374
rect 47248 37210 47448 39090
rect 47186 37200 47506 37210
rect 47186 36800 47198 37200
rect 47498 36800 47506 37200
rect 47186 36790 47506 36800
rect 47964 35752 48364 39990
rect 47964 35368 47974 35752
rect 48358 35368 48364 35752
rect 47248 32588 47448 34468
rect 47186 32578 47506 32588
rect 47186 32178 47198 32578
rect 47498 32178 47506 32578
rect 47186 32168 47506 32178
rect 47964 31130 48364 35368
rect 47964 30746 47974 31130
rect 48358 30746 48364 31130
rect 47248 27966 47448 29846
rect 47186 27956 47506 27966
rect 47186 27556 47198 27956
rect 47498 27556 47506 27956
rect 47186 27546 47506 27556
rect 44792 26124 44802 26508
rect 45186 26124 45192 26508
rect 44792 21886 45192 26124
rect 47964 26508 48364 30746
rect 47964 26124 47974 26508
rect 48358 26124 48364 26508
rect 47248 23344 47448 25224
rect 47186 23334 47506 23344
rect 47186 22934 47198 23334
rect 47498 22934 47506 23334
rect 47186 22924 47506 22934
rect 44792 21502 44802 21886
rect 45186 21502 45192 21886
rect 44792 17264 45192 21502
rect 47964 21886 48364 26124
rect 47964 21502 47974 21886
rect 48358 21502 48364 21886
rect 47248 18722 47448 20602
rect 47186 18712 47506 18722
rect 47186 18312 47198 18712
rect 47498 18312 47506 18712
rect 47186 18302 47506 18312
rect 44792 16880 44802 17264
rect 45186 16880 45192 17264
rect 44792 7420 45192 16880
rect 47964 17264 48364 21502
rect 48684 32570 49084 32590
rect 48684 32190 48700 32570
rect 49070 32190 49084 32570
rect 48684 18110 49084 32190
rect 51020 22750 51220 25224
rect 50958 22740 51278 22750
rect 50958 22340 50970 22740
rect 51270 22340 51278 22740
rect 50958 22330 51278 22340
rect 51020 18128 51220 20602
rect 48684 17730 48700 18110
rect 49070 17730 49084 18110
rect 48684 17720 49084 17730
rect 50958 18118 51278 18128
rect 50958 17718 50970 18118
rect 51270 17718 51278 18118
rect 50958 17708 51278 17718
rect 47964 16880 47974 17264
rect 48358 16880 48364 17264
rect 47248 14100 47448 15980
rect 47186 14090 47506 14100
rect 47186 13690 47198 14090
rect 47498 13690 47506 14090
rect 47186 13680 47506 13690
rect 47964 8050 48364 16880
rect 51020 13506 51220 15980
rect 50958 13496 51278 13506
rect 50958 13096 50970 13496
rect 51270 13096 51278 13496
rect 50958 13086 51278 13096
rect 47964 7670 47980 8050
rect 48350 7670 48364 8050
rect 47964 7660 48364 7670
rect 50650 12650 50890 12660
rect 50650 12260 51210 12650
rect 44790 7410 45192 7420
rect 44790 7030 44800 7410
rect 45180 7030 45192 7410
rect 44790 7020 45192 7030
rect 40420 5560 40430 5940
rect 40810 5560 40820 5940
rect 44190 6190 44592 6200
rect 44190 5810 44200 6190
rect 44580 5810 44592 6190
rect 44190 5800 44592 5810
rect 44792 5800 45192 7020
rect 46170 6790 46440 6800
rect 46170 6410 46180 6790
rect 46430 6410 46440 6790
rect 46170 6400 46440 6410
rect 40420 5550 40820 5560
rect 50650 5680 50890 12260
rect 38620 5410 38870 5420
rect 37410 4870 37420 5250
rect 37790 4870 37800 5250
rect 37410 4860 37800 4870
rect 50650 5390 50660 5680
rect 50880 5390 50890 5680
rect 36640 4340 36650 4720
rect 37040 4340 37050 4720
rect 36640 3470 37050 4340
rect 38310 3700 38540 4300
rect 38300 3690 38550 3700
rect 38300 3310 38310 3690
rect 38540 3310 38550 3690
rect 38300 3300 38550 3310
rect 46170 3640 46410 4280
rect 50650 4210 50890 5390
rect 50650 3830 50660 4210
rect 50880 3830 50890 4210
rect 50650 3820 50890 3830
rect 51000 4460 51240 11380
rect 51000 4070 51010 4460
rect 51230 4070 51240 4460
rect 46170 3630 46620 3640
rect 32870 2610 32880 2990
rect 33270 2610 33280 2990
rect 32870 2600 33280 2610
rect 27660 2540 28660 2550
rect 27660 2060 27670 2540
rect 28650 2060 28660 2540
rect 38310 2480 38540 3300
rect 46170 3250 46180 3630
rect 46610 3250 46620 3630
rect 46170 3240 46620 3250
rect 46170 3220 46410 3240
rect 38300 2470 38550 2480
rect 38300 2090 38310 2470
rect 38540 2090 38550 2470
rect 38300 2080 38550 2090
rect 27660 2050 28660 2060
rect 51000 1380 51240 4070
rect 50980 1370 51260 1380
rect 18200 1170 19200 1180
rect 1590 1150 2590 1160
rect 1590 670 1600 1150
rect 2580 670 2590 1150
rect 18200 690 18210 1170
rect 19190 690 19200 1170
rect 50980 1110 50990 1370
rect 51250 1110 51260 1370
rect 50980 1100 51260 1110
rect 51350 930 51410 40666
rect 51736 40374 52136 40600
rect 51736 39990 51746 40374
rect 52130 39990 52136 40374
rect 51736 35752 52136 39990
rect 51736 35368 51746 35752
rect 52130 35368 52136 35752
rect 51736 31130 52136 35368
rect 51736 30746 51746 31130
rect 52130 30746 52136 31130
rect 51736 6200 52136 30746
rect 52336 26508 52736 40600
rect 55508 40374 55908 40600
rect 55508 39990 55518 40374
rect 55902 39990 55908 40374
rect 52336 26124 52346 26508
rect 52730 26124 52736 26508
rect 52336 21886 52736 26124
rect 52336 21502 52346 21886
rect 52730 21502 52736 21886
rect 52336 17264 52736 21502
rect 52336 16880 52346 17264
rect 52730 16880 52736 17264
rect 52336 7620 52736 16880
rect 55508 35752 55908 39990
rect 59280 40374 59680 40600
rect 59280 39990 59290 40374
rect 59674 39990 59680 40374
rect 55508 35368 55518 35752
rect 55902 35368 55908 35752
rect 55508 31130 55908 35368
rect 55508 30746 55518 31130
rect 55902 30746 55908 31130
rect 55508 26508 55908 30746
rect 59280 35752 59680 39990
rect 63052 40374 63452 40600
rect 63052 39990 63062 40374
rect 63446 39990 63452 40374
rect 62336 37210 62536 39090
rect 62274 37200 62594 37210
rect 62274 36800 62286 37200
rect 62586 36800 62594 37200
rect 62274 36790 62594 36800
rect 59280 35368 59290 35752
rect 59674 35368 59680 35752
rect 59280 31130 59680 35368
rect 63052 35752 63452 39990
rect 66824 40374 67224 40600
rect 66824 39990 66834 40374
rect 67218 39990 67224 40374
rect 66108 37210 66308 39090
rect 66046 37200 66366 37210
rect 66046 36800 66058 37200
rect 66358 36800 66366 37200
rect 66046 36790 66366 36800
rect 63052 35368 63062 35752
rect 63446 35368 63452 35752
rect 62336 32588 62536 34468
rect 62274 32578 62594 32588
rect 62274 32178 62286 32578
rect 62586 32178 62594 32578
rect 62274 32168 62594 32178
rect 59280 30746 59290 31130
rect 59674 30746 59680 31130
rect 55508 26124 55518 26508
rect 55902 26124 55908 26508
rect 55508 21886 55908 26124
rect 55508 21502 55518 21886
rect 55902 21502 55908 21886
rect 55508 17264 55908 21502
rect 55508 16880 55518 17264
rect 55902 16880 55908 17264
rect 55508 16710 55908 16880
rect 56228 27940 56628 27970
rect 56228 27570 56240 27940
rect 56620 27570 56628 27940
rect 55508 16000 55910 16710
rect 51730 6190 52136 6200
rect 52330 7610 52736 7620
rect 52330 7230 52340 7610
rect 52720 7410 52736 7610
rect 52720 7230 52730 7410
rect 51730 5810 51740 6190
rect 52120 5810 52130 6190
rect 51730 5800 52130 5810
rect 52330 5800 52730 7230
rect 55510 5740 55910 16000
rect 56228 13480 56628 27570
rect 56228 13110 56240 13480
rect 56610 13110 56628 13480
rect 56228 13090 56628 13110
rect 59280 26508 59680 30746
rect 63052 31130 63452 35368
rect 66824 35752 67224 39990
rect 70596 40374 70996 40600
rect 70596 39990 70606 40374
rect 70990 39990 70996 40374
rect 66824 35368 66834 35752
rect 67218 35368 67224 35752
rect 66108 32588 66308 34468
rect 66046 32578 66366 32588
rect 66046 32178 66058 32578
rect 66358 32178 66366 32578
rect 66046 32168 66366 32178
rect 63052 30746 63062 31130
rect 63446 30746 63452 31130
rect 62336 27966 62536 29846
rect 62274 27956 62594 27966
rect 62274 27556 62286 27956
rect 62586 27556 62594 27956
rect 62274 27546 62594 27556
rect 59280 26124 59290 26508
rect 59674 26124 59680 26508
rect 59280 21886 59680 26124
rect 63052 26508 63452 30746
rect 66824 31130 67224 35368
rect 66824 30746 66834 31130
rect 67218 30746 67224 31130
rect 66108 27966 66308 29846
rect 66046 27956 66366 27966
rect 66046 27556 66058 27956
rect 66358 27556 66366 27956
rect 66046 27546 66366 27556
rect 63052 26124 63062 26508
rect 63446 26124 63452 26508
rect 62336 23344 62536 25224
rect 62274 23334 62594 23344
rect 62274 22934 62286 23334
rect 62586 22934 62594 23334
rect 62274 22924 62594 22934
rect 59280 21502 59290 21886
rect 59674 21502 59680 21886
rect 59280 17264 59680 21502
rect 63052 21886 63452 26124
rect 66824 26508 67224 30746
rect 66824 26124 66834 26508
rect 67218 26124 67224 26508
rect 66108 23344 66308 25224
rect 66046 23334 66366 23344
rect 66046 22934 66058 23334
rect 66358 22934 66366 23334
rect 66046 22924 66366 22934
rect 63052 21502 63062 21886
rect 63446 21502 63452 21886
rect 62336 18722 62536 20602
rect 62274 18712 62594 18722
rect 62274 18312 62286 18712
rect 62586 18312 62594 18712
rect 62274 18302 62594 18312
rect 63052 17800 63452 21502
rect 66824 21886 67224 26124
rect 70596 35752 70996 39990
rect 70596 35368 70606 35752
rect 70990 35368 70996 35752
rect 70596 31130 70996 35368
rect 70596 30746 70606 31130
rect 70990 30746 70996 31130
rect 69880 22750 70080 25224
rect 69818 22740 70138 22750
rect 69818 22340 69830 22740
rect 70130 22340 70138 22740
rect 69818 22330 70138 22340
rect 66824 21502 66834 21886
rect 67218 21502 67224 21886
rect 66108 18722 66308 20602
rect 66046 18712 66366 18722
rect 66046 18312 66058 18712
rect 66358 18312 66366 18712
rect 66046 18302 66366 18312
rect 59280 16880 59290 17264
rect 59674 16880 59680 17264
rect 55510 5390 55520 5740
rect 55900 5390 55910 5740
rect 55510 5340 55910 5390
rect 59280 10940 59680 16880
rect 63050 17264 63452 17800
rect 63050 16880 63062 17264
rect 63446 16880 63452 17264
rect 63050 16000 63452 16880
rect 66824 17264 67224 21502
rect 69880 18128 70080 20602
rect 69818 18118 70138 18128
rect 69818 17718 69830 18118
rect 70130 17718 70138 18118
rect 69818 17708 70138 17718
rect 66824 16880 66834 17264
rect 67218 16880 67224 17264
rect 66824 16000 67224 16880
rect 70596 16000 70996 30746
rect 71196 26508 71596 40600
rect 74368 40374 74768 40600
rect 74368 39990 74378 40374
rect 74762 39990 74768 40374
rect 71196 26124 71206 26508
rect 71590 26124 71596 26508
rect 71196 21886 71596 26124
rect 71196 21502 71206 21886
rect 71590 21502 71596 21886
rect 71196 17264 71596 21502
rect 71196 16880 71206 17264
rect 71590 16880 71596 17264
rect 71196 16000 71596 16880
rect 74368 35752 74768 39990
rect 78140 40374 78540 40600
rect 78140 39990 78150 40374
rect 78534 39990 78540 40374
rect 74368 35368 74378 35752
rect 74762 35368 74768 35752
rect 74368 31130 74768 35368
rect 74368 30746 74378 31130
rect 74762 30746 74768 31130
rect 74368 26508 74768 30746
rect 74368 26124 74378 26508
rect 74762 26124 74768 26508
rect 74368 21886 74768 26124
rect 78140 35752 78540 39990
rect 81912 40374 82312 40600
rect 81912 39990 81922 40374
rect 82306 39990 82312 40374
rect 78140 35368 78150 35752
rect 78534 35368 78540 35752
rect 78140 31130 78540 35368
rect 78140 30746 78150 31130
rect 78534 30746 78540 31130
rect 78140 26508 78540 30746
rect 78140 26124 78150 26508
rect 78534 26124 78540 26508
rect 75120 23370 75528 23380
rect 75120 22390 75130 23370
rect 75520 22390 75528 23370
rect 75120 22380 75528 22390
rect 74368 21502 74378 21886
rect 74762 21502 74768 21886
rect 74368 17264 74768 21502
rect 74368 16880 74378 17264
rect 74762 16880 74768 17264
rect 74368 16000 74768 16880
rect 62336 14100 62536 15980
rect 62274 14090 62594 14100
rect 62274 13690 62286 14090
rect 62586 13690 62594 14090
rect 62274 13680 62594 13690
rect 59280 10560 59290 10940
rect 59670 10560 59680 10940
rect 59280 6320 59680 10560
rect 59280 5930 59290 6320
rect 59670 5930 59680 6320
rect 53070 1020 53310 4360
rect 51780 1010 53310 1020
rect 51350 920 51600 930
rect 51350 710 51360 920
rect 51590 710 51600 920
rect 51780 850 51790 1010
rect 52040 850 53310 1010
rect 51780 840 53310 850
rect 51350 700 51600 710
rect 18200 680 19200 690
rect 1590 660 2590 670
rect 11340 490 12340 500
rect 7180 390 8780 400
rect 186 0 366 200
rect 4050 0 4230 200
rect 7180 10 7190 390
rect 8770 10 8780 390
rect 7180 0 8780 10
rect 11340 10 11350 490
rect 12330 10 12340 490
rect 11340 0 12340 10
rect 15240 490 16240 500
rect 15240 10 15250 490
rect 16230 10 16240 490
rect 15240 0 16240 10
rect 19460 490 20460 500
rect 19460 10 19470 490
rect 20450 10 20460 490
rect 19460 0 20460 10
rect 22960 490 23960 500
rect 22960 10 22970 490
rect 23950 10 23960 490
rect 22960 0 23960 10
rect 26820 490 27820 500
rect 26820 10 26830 490
rect 27810 10 27820 490
rect 53070 340 53310 840
rect 53390 1030 53630 4120
rect 53390 840 53400 1030
rect 53620 840 53630 1030
rect 53390 660 53630 840
rect 53720 980 53960 4400
rect 59280 3500 59680 5930
rect 63050 10940 63450 16000
rect 66108 14100 66308 15980
rect 66046 14090 66366 14100
rect 66046 13690 66058 14090
rect 66358 13690 66366 14090
rect 66046 13680 66366 13690
rect 66830 11430 67220 16000
rect 69880 13506 70080 15980
rect 69818 13496 70138 13506
rect 69818 13096 69830 13496
rect 70130 13096 70138 13496
rect 69818 13086 70138 13096
rect 66830 11050 66840 11430
rect 67210 11050 67220 11430
rect 66830 11040 67220 11050
rect 70600 12960 70990 16000
rect 70600 12770 70610 12960
rect 70980 12770 70990 12960
rect 63050 10560 63060 10940
rect 63440 10560 63450 10940
rect 63050 8480 63450 10560
rect 70600 10130 70990 12770
rect 70600 9940 70610 10130
rect 70980 9940 70990 10130
rect 70600 9650 70990 9940
rect 71200 12690 71590 16000
rect 71200 12500 71210 12690
rect 71580 12500 71590 12690
rect 71200 9860 71590 12500
rect 74370 10410 74760 16000
rect 74370 10020 74380 10410
rect 74750 10020 74760 10410
rect 74370 10010 74760 10020
rect 71200 9670 71210 9860
rect 71580 9670 71590 9860
rect 71200 9650 71590 9670
rect 63050 8160 63060 8480
rect 63440 8160 63450 8480
rect 63050 6320 63450 8160
rect 63050 5930 63060 6320
rect 63440 5930 63450 6320
rect 63050 4190 63450 5930
rect 59280 2860 59300 3500
rect 59660 2860 59680 3500
rect 65030 3810 65270 4140
rect 65030 3800 65490 3810
rect 65030 3220 65040 3800
rect 65480 3220 65490 3800
rect 65030 3210 65490 3220
rect 59280 2840 59680 2860
rect 75128 2180 75528 22380
rect 78140 21886 78540 26124
rect 78140 21502 78150 21886
rect 78534 21502 78540 21886
rect 78140 17264 78540 21502
rect 81912 35752 82312 39990
rect 85684 40374 86084 40600
rect 85684 39990 85694 40374
rect 86078 39990 86084 40374
rect 81912 35368 81922 35752
rect 82306 35368 82312 35752
rect 81912 31130 82312 35368
rect 81912 30746 81922 31130
rect 82306 30746 82312 31130
rect 81912 26508 82312 30746
rect 81912 26124 81922 26508
rect 82306 26124 82312 26508
rect 81912 21886 82312 26124
rect 81912 21502 81922 21886
rect 82306 21502 82312 21886
rect 78140 16880 78150 17264
rect 78534 16880 78540 17264
rect 78140 10940 78540 16880
rect 78140 10560 78150 10940
rect 78530 10560 78540 10940
rect 78140 5550 78540 10560
rect 78140 5210 78150 5550
rect 78530 5210 78540 5550
rect 78140 5200 78540 5210
rect 78900 18740 79300 18750
rect 78900 17760 78910 18740
rect 79290 17760 79300 18740
rect 75020 2170 75620 2180
rect 54290 1630 59850 1640
rect 54290 1420 54300 1630
rect 54540 1420 59360 1630
rect 59840 1420 59850 1630
rect 75020 1590 75030 2170
rect 75610 1590 75620 2170
rect 75020 1580 75620 1590
rect 54290 1410 59850 1420
rect 78900 1380 79300 17760
rect 81912 17264 82312 21502
rect 81912 16880 81922 17264
rect 82306 16880 82312 17264
rect 81912 8590 82312 16880
rect 85684 35752 86084 39990
rect 89456 40374 89856 40600
rect 89456 39990 89466 40374
rect 89850 39990 89856 40374
rect 88740 37210 88940 39090
rect 88678 37200 88998 37210
rect 88678 36800 88690 37200
rect 88990 36800 88998 37200
rect 88678 36790 88998 36800
rect 85684 35368 85694 35752
rect 86078 35368 86084 35752
rect 85684 31130 86084 35368
rect 89456 35752 89856 39990
rect 93228 40374 93628 40600
rect 93228 39990 93238 40374
rect 93622 39990 93628 40374
rect 92512 37210 92712 39090
rect 92450 37200 92770 37210
rect 92450 36800 92462 37200
rect 92762 36800 92770 37200
rect 92450 36790 92770 36800
rect 89456 35368 89466 35752
rect 89850 35368 89856 35752
rect 88740 32588 88940 34468
rect 88678 32578 88998 32588
rect 88678 32178 88690 32578
rect 88990 32178 88998 32578
rect 88678 32168 88998 32178
rect 85684 30746 85694 31130
rect 86078 30746 86084 31130
rect 85684 26508 86084 30746
rect 89456 31130 89856 35368
rect 93228 35752 93628 39990
rect 97000 40374 97400 40600
rect 97000 39990 97010 40374
rect 97394 39990 97400 40374
rect 96284 37210 96484 39090
rect 96222 37200 96542 37210
rect 96222 36800 96234 37200
rect 96534 36800 96542 37200
rect 96222 36790 96542 36800
rect 93228 35368 93238 35752
rect 93622 35368 93628 35752
rect 92512 32588 92712 34468
rect 92450 32578 92770 32588
rect 92450 32178 92462 32578
rect 92762 32178 92770 32578
rect 92450 32168 92770 32178
rect 89456 30746 89466 31130
rect 89850 30746 89856 31130
rect 88740 27966 88940 29846
rect 88678 27956 88998 27966
rect 88678 27556 88690 27956
rect 88990 27556 88998 27956
rect 88678 27546 88998 27556
rect 85684 26124 85694 26508
rect 86078 26124 86084 26508
rect 85684 21886 86084 26124
rect 89456 26508 89856 30746
rect 93228 31130 93628 35368
rect 97000 35752 97400 39990
rect 97000 35368 97010 35752
rect 97394 35368 97400 35752
rect 96284 32588 96484 34468
rect 96222 32578 96542 32588
rect 96222 32178 96234 32578
rect 96534 32178 96542 32578
rect 96222 32168 96542 32178
rect 93228 30746 93238 31130
rect 93622 30746 93628 31130
rect 92512 27966 92712 29846
rect 92450 27956 92770 27966
rect 92450 27556 92462 27956
rect 92762 27556 92770 27956
rect 92450 27546 92770 27556
rect 89456 26124 89466 26508
rect 89850 26124 89856 26508
rect 88740 23344 88940 25224
rect 88678 23334 88998 23344
rect 88678 22934 88690 23334
rect 88990 22934 88998 23334
rect 88678 22924 88998 22934
rect 85684 21502 85694 21886
rect 86078 21502 86084 21886
rect 85684 17264 86084 21502
rect 89456 21886 89856 26124
rect 93228 26508 93628 30746
rect 97000 31130 97400 35368
rect 97000 30746 97010 31130
rect 97394 30746 97400 31130
rect 96284 27966 96484 29846
rect 96222 27956 96542 27966
rect 96222 27556 96234 27956
rect 96534 27556 96542 27956
rect 96222 27546 96542 27556
rect 93228 26124 93238 26508
rect 93622 26124 93628 26508
rect 90130 24150 90660 24160
rect 90130 23470 90140 24150
rect 90650 23470 90660 24150
rect 90130 23460 90660 23470
rect 89456 21502 89466 21886
rect 89850 21502 89856 21886
rect 88740 18722 88940 20602
rect 88678 18712 88998 18722
rect 88678 18312 88690 18712
rect 88990 18312 88998 18712
rect 88678 18302 88998 18312
rect 85684 16880 85694 17264
rect 86078 16880 86084 17264
rect 81912 8350 81920 8590
rect 82300 8350 82312 8590
rect 81912 8340 82312 8350
rect 82670 14090 83070 15960
rect 82670 13110 82680 14090
rect 83060 13700 83070 14090
rect 83060 13110 83072 13700
rect 80120 6490 81380 6730
rect 82670 2020 83072 13110
rect 85684 12640 86084 16880
rect 89456 17264 89856 21502
rect 89456 16880 89466 17264
rect 89850 16880 89856 17264
rect 88740 14100 88940 15980
rect 88678 14090 88998 14100
rect 88678 13690 88690 14090
rect 88990 13690 88998 14090
rect 88678 13680 88998 13690
rect 85684 12270 85700 12640
rect 86070 12270 86084 12640
rect 85684 6580 86084 12270
rect 89456 12640 89856 16880
rect 89456 12270 89470 12640
rect 89840 12270 89856 12640
rect 85684 6190 85690 6580
rect 86070 6190 86084 6580
rect 85684 6180 86084 6190
rect 86520 9340 86890 9350
rect 86520 8960 86530 9340
rect 86880 8960 86890 9340
rect 86520 4960 86890 8960
rect 86520 4590 86530 4960
rect 86880 4590 86890 4960
rect 86520 4580 86890 4590
rect 88580 2180 89020 6760
rect 89456 3260 89856 12270
rect 90216 8020 90616 23460
rect 92512 23344 92712 25224
rect 92450 23334 92770 23344
rect 92450 22934 92462 23334
rect 92762 22934 92770 23334
rect 92450 22924 92770 22934
rect 93228 21886 93628 26124
rect 97000 26508 97400 30746
rect 97000 26124 97010 26508
rect 97394 26124 97400 26508
rect 96284 23344 96484 25224
rect 96222 23334 96542 23344
rect 96222 22934 96234 23334
rect 96534 22934 96542 23334
rect 96222 22924 96542 22934
rect 93228 21502 93238 21886
rect 93622 21502 93628 21886
rect 92512 18722 92712 20602
rect 92450 18712 92770 18722
rect 92450 18312 92462 18712
rect 92762 18312 92770 18712
rect 92450 18302 92770 18312
rect 93228 17264 93628 21502
rect 97000 21886 97400 26124
rect 97000 21502 97010 21886
rect 97394 21502 97400 21886
rect 93900 19520 94430 19530
rect 93900 18840 93910 19520
rect 94420 18840 94430 19520
rect 93900 18830 94430 18840
rect 93228 16880 93238 17264
rect 93622 16880 93628 17264
rect 92512 14100 92712 15980
rect 92450 14090 92770 14100
rect 92450 13690 92462 14090
rect 92762 13690 92770 14090
rect 92450 13680 92770 13690
rect 90216 7300 90220 8020
rect 90600 7300 90616 8020
rect 90216 7290 90616 7300
rect 89456 2870 89470 3260
rect 89840 2870 89856 3260
rect 89456 2860 89856 2870
rect 88500 2170 89100 2180
rect 78800 1370 79400 1380
rect 53720 740 54560 980
rect 78800 790 78810 1370
rect 79390 790 79400 1370
rect 78800 780 79400 790
rect 82670 680 83070 2020
rect 88500 1590 88510 2170
rect 89090 1590 89100 2170
rect 88500 1580 89100 1590
rect 92320 1390 92760 6760
rect 93228 3260 93628 16880
rect 93988 8020 94388 18830
rect 96284 18722 96484 20602
rect 96222 18712 96542 18722
rect 96222 18312 96234 18712
rect 96534 18312 96542 18712
rect 96222 18302 96542 18312
rect 97000 17264 97400 21502
rect 97000 16880 97010 17264
rect 97394 16880 97400 17264
rect 96284 14100 96484 15980
rect 96222 14090 96542 14100
rect 96222 13690 96234 14090
rect 96534 13690 96542 14090
rect 96222 13680 96542 13690
rect 93988 7300 94000 8020
rect 94380 7300 94388 8020
rect 93988 7290 94388 7300
rect 97000 10940 97400 16880
rect 97000 10560 97010 10940
rect 97390 10560 97400 10940
rect 93228 2870 93240 3260
rect 93620 2870 93628 3260
rect 93228 2860 93628 2870
rect 92240 1380 92840 1390
rect 92240 800 92250 1380
rect 92830 800 92840 1380
rect 92240 790 92840 800
rect 96140 690 96580 6760
rect 97000 3930 97400 10560
rect 97760 14680 98160 14700
rect 97760 13700 97770 14680
rect 98150 13700 98160 14680
rect 97760 8020 98160 13700
rect 97760 7300 97770 8020
rect 98150 7300 98160 8020
rect 97760 7290 98160 7300
rect 97000 3530 97010 3930
rect 97390 3530 97400 3930
rect 97000 3520 97400 3530
rect 96060 680 96660 690
rect 82570 670 83170 680
rect 53390 420 54490 660
rect 53070 110 54650 340
rect 82570 90 82580 670
rect 83160 90 83170 670
rect 96060 100 96070 680
rect 96650 100 96660 680
rect 96060 90 96660 100
rect 82570 80 83170 90
rect 26820 0 27820 10
use mosbius_col6  mosbius_col6_2
timestamp 1757289701
transform 1 0 64370 0 1 36332
box -146 -32354 3794 8020
use mosbius_col6  mosbius_col6_3
timestamp 1757289701
transform 1 0 68142 0 1 36332
box -146 -32354 3794 8020
use mosbius_col7  mosbius_col7_9
timestamp 1757297520
transform 1 0 7790 0 1 36332
box -146 -32354 3794 8020
use mosbius_col7  mosbius_col7_10
timestamp 1757297520
transform 1 0 11562 0 1 36332
box -146 -32354 3794 8020
use mosbius_col7  mosbius_col7_11
timestamp 1757297520
transform 1 0 37966 0 1 36332
box -146 -32354 3794 8020
use mosbius_col7  mosbius_col7_12
timestamp 1757297520
transform 1 0 45510 0 1 36332
box -146 -32354 3794 8020
use mosbius_col7  mosbius_col7_13
timestamp 1757297520
transform 1 0 41738 0 1 36332
box -146 -32354 3794 8020
use mosbius_col7  mosbius_col7_14
timestamp 1757297520
transform 1 0 49282 0 1 36332
box -146 -32354 3794 8020
use mosbius_col7  mosbius_col7_15
timestamp 1757297520
transform 1 0 71914 0 1 36332
box -146 -32354 3794 8020
use mosbius_col7  mosbius_col7_16
timestamp 1757297520
transform 1 0 83230 0 1 36332
box -146 -32354 3794 8020
use mosbius_col8  mosbius_col8_3
timestamp 1757297674
transform 1 0 246 0 1 36332
box -146 -32354 3794 8020
use mosbius_col8  mosbius_col8_4
timestamp 1757297674
transform 1 0 4018 0 1 36332
box -146 -32354 3794 8020
use mosbius_col8  mosbius_col8_11
timestamp 1757297674
transform 1 0 15334 0 1 36332
box -146 -32354 3794 8020
use mosbius_col8  mosbius_col8_12
timestamp 1757297674
transform 1 0 30422 0 1 36332
box -146 -32354 3794 8020
use mosbius_col8  mosbius_col8_13
timestamp 1757297674
transform 1 0 26650 0 1 36332
box -146 -32354 3794 8020
use mosbius_col8  mosbius_col8_14
timestamp 1757297674
transform 1 0 22878 0 1 36332
box -146 -32354 3794 8020
use mosbius_col8  mosbius_col8_18
timestamp 1757297674
transform 1 0 19106 0 1 36332
box -146 -32354 3794 8020
use mosbius_col8  mosbius_col8_19
timestamp 1757297674
transform 1 0 34194 0 1 36332
box -146 -32354 3794 8020
use mosbius_col8  mosbius_col8_20
timestamp 1757297674
transform 1 0 60598 0 1 36332
box -146 -32354 3794 8020
use mosbius_col8  mosbius_col8_21
timestamp 1757297674
transform 1 0 56826 0 1 36332
box -146 -32354 3794 8020
use mosbius_col8  mosbius_col8_24
timestamp 1757297674
transform 1 0 53054 0 1 36332
box -146 -32354 3794 8020
use mosbius_col8  mosbius_col8_26
timestamp 1757297674
transform 1 0 75686 0 1 36332
box -146 -32354 3794 8020
use mosbius_col8  mosbius_col8_27
timestamp 1757297674
transform 1 0 79458 0 1 36332
box -146 -32354 3794 8020
use mosbius_col8  mosbius_col8_28
timestamp 1757297674
transform 1 0 90774 0 1 36332
box -146 -32354 3794 8020
use mosbius_col8  mosbius_col8_29
timestamp 1757297674
transform 1 0 94546 0 1 36332
box -146 -32354 3794 8020
use mosbius_col8  mosbius_col8_30
timestamp 1757297674
transform 1 0 87002 0 1 36332
box -146 -32354 3794 8020
use sky130_fd_pr__nfet_01v8_EDB9KC  sky130_fd_pr__nfet_01v8_EDB9KC_0
timestamp 1757297086
transform 1 0 52538 0 1 929
box -211 -252 211 252
use sky130_fd_pr__nfet_g5v0d10v5_8ML6AG  sky130_fd_pr__nfet_g5v0d10v5_8ML6AG_2
timestamp 1757283562
transform 1 0 40671 0 1 6608
box -1621 -758 1621 758
use sky130_fd_pr__nfet_g5v0d10v5_8ML6AG  sky130_fd_pr__nfet_g5v0d10v5_8ML6AG_3
timestamp 1757283562
transform 1 0 49071 0 1 6608
box -1621 -758 1621 758
use sky130_fd_pr__nfet_g5v0d10v5_8263FJ  sky130_fd_pr__nfet_g5v0d10v5_8263FJ_1
timestamp 1757283562
transform -1 0 9573 0 -1 5967
box -673 -1367 673 1367
use sky130_fd_pr__nfet_g5v0d10v5_8263FJ  sky130_fd_pr__nfet_g5v0d10v5_8263FJ_3
timestamp 1757283562
transform -1 0 13273 0 -1 5967
box -673 -1367 673 1367
use sky130_fd_pr__nfet_g5v0d10v5_CLGMFJ  sky130_fd_pr__nfet_g5v0d10v5_CLGMFJ_1
timestamp 1757283562
transform 1 0 42411 0 1 3167
box -3811 -1367 3811 1367
use sky130_fd_pr__pfet_01v8_hvt_UAQRRG  sky130_fd_pr__pfet_01v8_hvt_UAQRRG_0
timestamp 1757297086
transform 1 0 52081 0 1 929
box -211 -319 211 319
use sky130_fd_pr__pfet_g5v0d10v5_AA5R3U  sky130_fd_pr__pfet_g5v0d10v5_AA5R3U_2
timestamp 1757283562
transform 1 0 68183 0 1 11315
box -2283 -1415 2283 1415
use sky130_fd_pr__pfet_g5v0d10v5_FGL9HY  sky130_fd_pr__pfet_g5v0d10v5_FGL9HY_0
timestamp 1757283562
transform 1 0 85223 0 1 6725
box -1335 -1415 1335 1415
use sky130_fd_pr__pfet_g5v0d10v5_FGL9HY  sky130_fd_pr__pfet_g5v0d10v5_FGL9HY_3
timestamp 1757283562
transform 1 0 85213 0 1 3405
box -1335 -1415 1335 1415
use sky130_fd_pr__pfet_g5v0d10v5_N4SDRF  sky130_fd_pr__pfet_g5v0d10v5_N4SDRF_1
timestamp 1757283562
transform -1 0 70241 0 -1 5551
box -3841 -2651 3841 2651
use sky130_fd_pr__pfet_g5v0d10v5_R4AJ4P  sky130_fd_pr__pfet_g5v0d10v5_R4AJ4P_1
timestamp 1757283562
transform 1 0 48735 0 1 3115
box -2035 -1415 2035 1415
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_0
timestamp 1757289622
transform -1 0 27002 0 -1 44706
box -38 -48 314 592
use tt_asw_3v3  tt_asw_3v3_0
timestamp 1757289622
transform 0 -1 58720 1 0 82
box 0 0 3612 4352
<< labels >>
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 620 43980 800 44160 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 940 43980 1120 44160 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
flabel metal4 300 43980 480 44160 1 FreeSans 400 0 0 0 VDPWR
port 54 nsew power bidirectional
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 98624 45152
<< end >>
