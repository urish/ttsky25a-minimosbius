magic
tech sky130A
magscale 1 2
timestamp 1757283562
<< pwell >>
rect -673 -1367 673 1367
<< mvnmos >>
rect -445 109 -345 1109
rect -287 109 -187 1109
rect -129 109 -29 1109
rect 29 109 129 1109
rect 187 109 287 1109
rect 345 109 445 1109
rect -445 -1109 -345 -109
rect -287 -1109 -187 -109
rect -129 -1109 -29 -109
rect 29 -1109 129 -109
rect 187 -1109 287 -109
rect 345 -1109 445 -109
<< mvndiff >>
rect -503 1097 -445 1109
rect -503 121 -491 1097
rect -457 121 -445 1097
rect -503 109 -445 121
rect -345 1097 -287 1109
rect -345 121 -333 1097
rect -299 121 -287 1097
rect -345 109 -287 121
rect -187 1097 -129 1109
rect -187 121 -175 1097
rect -141 121 -129 1097
rect -187 109 -129 121
rect -29 1097 29 1109
rect -29 121 -17 1097
rect 17 121 29 1097
rect -29 109 29 121
rect 129 1097 187 1109
rect 129 121 141 1097
rect 175 121 187 1097
rect 129 109 187 121
rect 287 1097 345 1109
rect 287 121 299 1097
rect 333 121 345 1097
rect 287 109 345 121
rect 445 1097 503 1109
rect 445 121 457 1097
rect 491 121 503 1097
rect 445 109 503 121
rect -503 -121 -445 -109
rect -503 -1097 -491 -121
rect -457 -1097 -445 -121
rect -503 -1109 -445 -1097
rect -345 -121 -287 -109
rect -345 -1097 -333 -121
rect -299 -1097 -287 -121
rect -345 -1109 -287 -1097
rect -187 -121 -129 -109
rect -187 -1097 -175 -121
rect -141 -1097 -129 -121
rect -187 -1109 -129 -1097
rect -29 -121 29 -109
rect -29 -1097 -17 -121
rect 17 -1097 29 -121
rect -29 -1109 29 -1097
rect 129 -121 187 -109
rect 129 -1097 141 -121
rect 175 -1097 187 -121
rect 129 -1109 187 -1097
rect 287 -121 345 -109
rect 287 -1097 299 -121
rect 333 -1097 345 -121
rect 287 -1109 345 -1097
rect 445 -121 503 -109
rect 445 -1097 457 -121
rect 491 -1097 503 -121
rect 445 -1109 503 -1097
<< mvndiffc >>
rect -491 121 -457 1097
rect -333 121 -299 1097
rect -175 121 -141 1097
rect -17 121 17 1097
rect 141 121 175 1097
rect 299 121 333 1097
rect 457 121 491 1097
rect -491 -1097 -457 -121
rect -333 -1097 -299 -121
rect -175 -1097 -141 -121
rect -17 -1097 17 -121
rect 141 -1097 175 -121
rect 299 -1097 333 -121
rect 457 -1097 491 -121
<< mvpsubdiff >>
rect -637 1319 637 1331
rect -637 1285 -529 1319
rect 529 1285 637 1319
rect -637 1273 637 1285
rect -637 1223 -579 1273
rect -637 -1223 -625 1223
rect -591 -1223 -579 1223
rect 579 1223 637 1273
rect -637 -1273 -579 -1223
rect 579 -1223 591 1223
rect 625 -1223 637 1223
rect 579 -1273 637 -1223
rect -637 -1285 637 -1273
rect -637 -1319 -529 -1285
rect 529 -1319 637 -1285
rect -637 -1331 637 -1319
<< mvpsubdiffcont >>
rect -529 1285 529 1319
rect -625 -1223 -591 1223
rect 591 -1223 625 1223
rect -529 -1319 529 -1285
<< poly >>
rect -445 1181 -345 1197
rect -445 1147 -429 1181
rect -361 1147 -345 1181
rect -445 1109 -345 1147
rect -287 1181 -187 1197
rect -287 1147 -271 1181
rect -203 1147 -187 1181
rect -287 1109 -187 1147
rect -129 1181 -29 1197
rect -129 1147 -113 1181
rect -45 1147 -29 1181
rect -129 1109 -29 1147
rect 29 1181 129 1197
rect 29 1147 45 1181
rect 113 1147 129 1181
rect 29 1109 129 1147
rect 187 1181 287 1197
rect 187 1147 203 1181
rect 271 1147 287 1181
rect 187 1109 287 1147
rect 345 1181 445 1197
rect 345 1147 361 1181
rect 429 1147 445 1181
rect 345 1109 445 1147
rect -445 71 -345 109
rect -445 37 -429 71
rect -361 37 -345 71
rect -445 21 -345 37
rect -287 71 -187 109
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 109
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 109
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 109
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect 345 71 445 109
rect 345 37 361 71
rect 429 37 445 71
rect 345 21 445 37
rect -445 -37 -345 -21
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -445 -109 -345 -71
rect -287 -37 -187 -21
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -287 -109 -187 -71
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -109 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -109 129 -71
rect 187 -37 287 -21
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 187 -109 287 -71
rect 345 -37 445 -21
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 345 -109 445 -71
rect -445 -1147 -345 -1109
rect -445 -1181 -429 -1147
rect -361 -1181 -345 -1147
rect -445 -1197 -345 -1181
rect -287 -1147 -187 -1109
rect -287 -1181 -271 -1147
rect -203 -1181 -187 -1147
rect -287 -1197 -187 -1181
rect -129 -1147 -29 -1109
rect -129 -1181 -113 -1147
rect -45 -1181 -29 -1147
rect -129 -1197 -29 -1181
rect 29 -1147 129 -1109
rect 29 -1181 45 -1147
rect 113 -1181 129 -1147
rect 29 -1197 129 -1181
rect 187 -1147 287 -1109
rect 187 -1181 203 -1147
rect 271 -1181 287 -1147
rect 187 -1197 287 -1181
rect 345 -1147 445 -1109
rect 345 -1181 361 -1147
rect 429 -1181 445 -1147
rect 345 -1197 445 -1181
<< polycont >>
rect -429 1147 -361 1181
rect -271 1147 -203 1181
rect -113 1147 -45 1181
rect 45 1147 113 1181
rect 203 1147 271 1181
rect 361 1147 429 1181
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect -429 -1181 -361 -1147
rect -271 -1181 -203 -1147
rect -113 -1181 -45 -1147
rect 45 -1181 113 -1147
rect 203 -1181 271 -1147
rect 361 -1181 429 -1147
<< locali >>
rect -625 1285 -529 1319
rect 529 1285 625 1319
rect -625 1223 -591 1285
rect 591 1223 625 1285
rect -445 1147 -429 1181
rect -361 1147 -345 1181
rect -287 1147 -271 1181
rect -203 1147 -187 1181
rect -129 1147 -113 1181
rect -45 1147 -29 1181
rect 29 1147 45 1181
rect 113 1147 129 1181
rect 187 1147 203 1181
rect 271 1147 287 1181
rect 345 1147 361 1181
rect 429 1147 445 1181
rect -491 1097 -457 1113
rect -491 105 -457 121
rect -333 1097 -299 1113
rect -333 105 -299 121
rect -175 1097 -141 1113
rect -175 105 -141 121
rect -17 1097 17 1113
rect -17 105 17 121
rect 141 1097 175 1113
rect 141 105 175 121
rect 299 1097 333 1113
rect 299 105 333 121
rect 457 1097 491 1113
rect 457 105 491 121
rect -445 37 -429 71
rect -361 37 -345 71
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect 345 37 361 71
rect 429 37 445 71
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 345 -71 361 -37
rect 429 -71 445 -37
rect -491 -121 -457 -105
rect -491 -1113 -457 -1097
rect -333 -121 -299 -105
rect -333 -1113 -299 -1097
rect -175 -121 -141 -105
rect -175 -1113 -141 -1097
rect -17 -121 17 -105
rect -17 -1113 17 -1097
rect 141 -121 175 -105
rect 141 -1113 175 -1097
rect 299 -121 333 -105
rect 299 -1113 333 -1097
rect 457 -121 491 -105
rect 457 -1113 491 -1097
rect -445 -1181 -429 -1147
rect -361 -1181 -345 -1147
rect -287 -1181 -271 -1147
rect -203 -1181 -187 -1147
rect -129 -1181 -113 -1147
rect -45 -1181 -29 -1147
rect 29 -1181 45 -1147
rect 113 -1181 129 -1147
rect 187 -1181 203 -1147
rect 271 -1181 287 -1147
rect 345 -1181 361 -1147
rect 429 -1181 445 -1147
rect -625 -1285 -591 -1223
rect 591 -1285 625 -1223
rect -625 -1319 -529 -1285
rect 529 -1319 625 -1285
<< viali >>
rect -429 1147 -361 1181
rect -271 1147 -203 1181
rect -113 1147 -45 1181
rect 45 1147 113 1181
rect 203 1147 271 1181
rect 361 1147 429 1181
rect -491 121 -457 1097
rect -333 121 -299 1097
rect -175 121 -141 1097
rect -17 121 17 1097
rect 141 121 175 1097
rect 299 121 333 1097
rect 457 121 491 1097
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect -491 -1097 -457 -121
rect -333 -1097 -299 -121
rect -175 -1097 -141 -121
rect -17 -1097 17 -121
rect 141 -1097 175 -121
rect 299 -1097 333 -121
rect 457 -1097 491 -121
rect -429 -1181 -361 -1147
rect -271 -1181 -203 -1147
rect -113 -1181 -45 -1147
rect 45 -1181 113 -1147
rect 203 -1181 271 -1147
rect 361 -1181 429 -1147
<< metal1 >>
rect -441 1181 -349 1187
rect -441 1147 -429 1181
rect -361 1147 -349 1181
rect -441 1141 -349 1147
rect -283 1181 -191 1187
rect -283 1147 -271 1181
rect -203 1147 -191 1181
rect -283 1141 -191 1147
rect -125 1181 -33 1187
rect -125 1147 -113 1181
rect -45 1147 -33 1181
rect -125 1141 -33 1147
rect 33 1181 125 1187
rect 33 1147 45 1181
rect 113 1147 125 1181
rect 33 1141 125 1147
rect 191 1181 283 1187
rect 191 1147 203 1181
rect 271 1147 283 1181
rect 191 1141 283 1147
rect 349 1181 441 1187
rect 349 1147 361 1181
rect 429 1147 441 1181
rect 349 1141 441 1147
rect -497 1097 -451 1109
rect -497 121 -491 1097
rect -457 121 -451 1097
rect -497 109 -451 121
rect -339 1097 -293 1109
rect -339 121 -333 1097
rect -299 121 -293 1097
rect -339 109 -293 121
rect -181 1097 -135 1109
rect -181 121 -175 1097
rect -141 121 -135 1097
rect -181 109 -135 121
rect -23 1097 23 1109
rect -23 121 -17 1097
rect 17 121 23 1097
rect -23 109 23 121
rect 135 1097 181 1109
rect 135 121 141 1097
rect 175 121 181 1097
rect 135 109 181 121
rect 293 1097 339 1109
rect 293 121 299 1097
rect 333 121 339 1097
rect 293 109 339 121
rect 451 1097 497 1109
rect 451 121 457 1097
rect 491 121 497 1097
rect 451 109 497 121
rect -441 71 -349 77
rect -441 37 -429 71
rect -361 37 -349 71
rect -441 31 -349 37
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect 349 71 441 77
rect 349 37 361 71
rect 429 37 441 71
rect 349 31 441 37
rect -441 -37 -349 -31
rect -441 -71 -429 -37
rect -361 -71 -349 -37
rect -441 -77 -349 -71
rect -283 -37 -191 -31
rect -283 -71 -271 -37
rect -203 -71 -191 -37
rect -283 -77 -191 -71
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect 191 -37 283 -31
rect 191 -71 203 -37
rect 271 -71 283 -37
rect 191 -77 283 -71
rect 349 -37 441 -31
rect 349 -71 361 -37
rect 429 -71 441 -37
rect 349 -77 441 -71
rect -497 -121 -451 -109
rect -497 -1097 -491 -121
rect -457 -1097 -451 -121
rect -497 -1109 -451 -1097
rect -339 -121 -293 -109
rect -339 -1097 -333 -121
rect -299 -1097 -293 -121
rect -339 -1109 -293 -1097
rect -181 -121 -135 -109
rect -181 -1097 -175 -121
rect -141 -1097 -135 -121
rect -181 -1109 -135 -1097
rect -23 -121 23 -109
rect -23 -1097 -17 -121
rect 17 -1097 23 -121
rect -23 -1109 23 -1097
rect 135 -121 181 -109
rect 135 -1097 141 -121
rect 175 -1097 181 -121
rect 135 -1109 181 -1097
rect 293 -121 339 -109
rect 293 -1097 299 -121
rect 333 -1097 339 -121
rect 293 -1109 339 -1097
rect 451 -121 497 -109
rect 451 -1097 457 -121
rect 491 -1097 497 -121
rect 451 -1109 497 -1097
rect -441 -1147 -349 -1141
rect -441 -1181 -429 -1147
rect -361 -1181 -349 -1147
rect -441 -1187 -349 -1181
rect -283 -1147 -191 -1141
rect -283 -1181 -271 -1147
rect -203 -1181 -191 -1147
rect -283 -1187 -191 -1181
rect -125 -1147 -33 -1141
rect -125 -1181 -113 -1147
rect -45 -1181 -33 -1147
rect -125 -1187 -33 -1181
rect 33 -1147 125 -1141
rect 33 -1181 45 -1147
rect 113 -1181 125 -1147
rect 33 -1187 125 -1181
rect 191 -1147 283 -1141
rect 191 -1181 203 -1147
rect 271 -1181 283 -1147
rect 191 -1187 283 -1181
rect 349 -1147 441 -1141
rect 349 -1181 361 -1147
rect 429 -1181 441 -1147
rect 349 -1187 441 -1181
<< properties >>
string FIXED_BBOX -608 -1302 608 1302
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.50 m 2 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
