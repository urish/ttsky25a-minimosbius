magic
tech sky130A
magscale 1 2
timestamp 1757051612
<< pwell >>
rect -1147 -1367 1147 1367
<< mvnmos >>
rect -919 109 -819 1109
rect -761 109 -661 1109
rect -603 109 -503 1109
rect -445 109 -345 1109
rect -287 109 -187 1109
rect -129 109 -29 1109
rect 29 109 129 1109
rect 187 109 287 1109
rect 345 109 445 1109
rect 503 109 603 1109
rect 661 109 761 1109
rect 819 109 919 1109
rect -919 -1109 -819 -109
rect -761 -1109 -661 -109
rect -603 -1109 -503 -109
rect -445 -1109 -345 -109
rect -287 -1109 -187 -109
rect -129 -1109 -29 -109
rect 29 -1109 129 -109
rect 187 -1109 287 -109
rect 345 -1109 445 -109
rect 503 -1109 603 -109
rect 661 -1109 761 -109
rect 819 -1109 919 -109
<< mvndiff >>
rect -977 1097 -919 1109
rect -977 121 -965 1097
rect -931 121 -919 1097
rect -977 109 -919 121
rect -819 1097 -761 1109
rect -819 121 -807 1097
rect -773 121 -761 1097
rect -819 109 -761 121
rect -661 1097 -603 1109
rect -661 121 -649 1097
rect -615 121 -603 1097
rect -661 109 -603 121
rect -503 1097 -445 1109
rect -503 121 -491 1097
rect -457 121 -445 1097
rect -503 109 -445 121
rect -345 1097 -287 1109
rect -345 121 -333 1097
rect -299 121 -287 1097
rect -345 109 -287 121
rect -187 1097 -129 1109
rect -187 121 -175 1097
rect -141 121 -129 1097
rect -187 109 -129 121
rect -29 1097 29 1109
rect -29 121 -17 1097
rect 17 121 29 1097
rect -29 109 29 121
rect 129 1097 187 1109
rect 129 121 141 1097
rect 175 121 187 1097
rect 129 109 187 121
rect 287 1097 345 1109
rect 287 121 299 1097
rect 333 121 345 1097
rect 287 109 345 121
rect 445 1097 503 1109
rect 445 121 457 1097
rect 491 121 503 1097
rect 445 109 503 121
rect 603 1097 661 1109
rect 603 121 615 1097
rect 649 121 661 1097
rect 603 109 661 121
rect 761 1097 819 1109
rect 761 121 773 1097
rect 807 121 819 1097
rect 761 109 819 121
rect 919 1097 977 1109
rect 919 121 931 1097
rect 965 121 977 1097
rect 919 109 977 121
rect -977 -121 -919 -109
rect -977 -1097 -965 -121
rect -931 -1097 -919 -121
rect -977 -1109 -919 -1097
rect -819 -121 -761 -109
rect -819 -1097 -807 -121
rect -773 -1097 -761 -121
rect -819 -1109 -761 -1097
rect -661 -121 -603 -109
rect -661 -1097 -649 -121
rect -615 -1097 -603 -121
rect -661 -1109 -603 -1097
rect -503 -121 -445 -109
rect -503 -1097 -491 -121
rect -457 -1097 -445 -121
rect -503 -1109 -445 -1097
rect -345 -121 -287 -109
rect -345 -1097 -333 -121
rect -299 -1097 -287 -121
rect -345 -1109 -287 -1097
rect -187 -121 -129 -109
rect -187 -1097 -175 -121
rect -141 -1097 -129 -121
rect -187 -1109 -129 -1097
rect -29 -121 29 -109
rect -29 -1097 -17 -121
rect 17 -1097 29 -121
rect -29 -1109 29 -1097
rect 129 -121 187 -109
rect 129 -1097 141 -121
rect 175 -1097 187 -121
rect 129 -1109 187 -1097
rect 287 -121 345 -109
rect 287 -1097 299 -121
rect 333 -1097 345 -121
rect 287 -1109 345 -1097
rect 445 -121 503 -109
rect 445 -1097 457 -121
rect 491 -1097 503 -121
rect 445 -1109 503 -1097
rect 603 -121 661 -109
rect 603 -1097 615 -121
rect 649 -1097 661 -121
rect 603 -1109 661 -1097
rect 761 -121 819 -109
rect 761 -1097 773 -121
rect 807 -1097 819 -121
rect 761 -1109 819 -1097
rect 919 -121 977 -109
rect 919 -1097 931 -121
rect 965 -1097 977 -121
rect 919 -1109 977 -1097
<< mvndiffc >>
rect -965 121 -931 1097
rect -807 121 -773 1097
rect -649 121 -615 1097
rect -491 121 -457 1097
rect -333 121 -299 1097
rect -175 121 -141 1097
rect -17 121 17 1097
rect 141 121 175 1097
rect 299 121 333 1097
rect 457 121 491 1097
rect 615 121 649 1097
rect 773 121 807 1097
rect 931 121 965 1097
rect -965 -1097 -931 -121
rect -807 -1097 -773 -121
rect -649 -1097 -615 -121
rect -491 -1097 -457 -121
rect -333 -1097 -299 -121
rect -175 -1097 -141 -121
rect -17 -1097 17 -121
rect 141 -1097 175 -121
rect 299 -1097 333 -121
rect 457 -1097 491 -121
rect 615 -1097 649 -121
rect 773 -1097 807 -121
rect 931 -1097 965 -121
<< mvpsubdiff >>
rect -1111 1319 1111 1331
rect -1111 1285 -1003 1319
rect 1003 1285 1111 1319
rect -1111 1273 1111 1285
rect -1111 1223 -1053 1273
rect -1111 -1223 -1099 1223
rect -1065 -1223 -1053 1223
rect 1053 1223 1111 1273
rect -1111 -1273 -1053 -1223
rect 1053 -1223 1065 1223
rect 1099 -1223 1111 1223
rect 1053 -1273 1111 -1223
rect -1111 -1285 1111 -1273
rect -1111 -1319 -1003 -1285
rect 1003 -1319 1111 -1285
rect -1111 -1331 1111 -1319
<< mvpsubdiffcont >>
rect -1003 1285 1003 1319
rect -1099 -1223 -1065 1223
rect 1065 -1223 1099 1223
rect -1003 -1319 1003 -1285
<< poly >>
rect -919 1181 -819 1197
rect -919 1147 -903 1181
rect -835 1147 -819 1181
rect -919 1109 -819 1147
rect -761 1181 -661 1197
rect -761 1147 -745 1181
rect -677 1147 -661 1181
rect -761 1109 -661 1147
rect -603 1181 -503 1197
rect -603 1147 -587 1181
rect -519 1147 -503 1181
rect -603 1109 -503 1147
rect -445 1181 -345 1197
rect -445 1147 -429 1181
rect -361 1147 -345 1181
rect -445 1109 -345 1147
rect -287 1181 -187 1197
rect -287 1147 -271 1181
rect -203 1147 -187 1181
rect -287 1109 -187 1147
rect -129 1181 -29 1197
rect -129 1147 -113 1181
rect -45 1147 -29 1181
rect -129 1109 -29 1147
rect 29 1181 129 1197
rect 29 1147 45 1181
rect 113 1147 129 1181
rect 29 1109 129 1147
rect 187 1181 287 1197
rect 187 1147 203 1181
rect 271 1147 287 1181
rect 187 1109 287 1147
rect 345 1181 445 1197
rect 345 1147 361 1181
rect 429 1147 445 1181
rect 345 1109 445 1147
rect 503 1181 603 1197
rect 503 1147 519 1181
rect 587 1147 603 1181
rect 503 1109 603 1147
rect 661 1181 761 1197
rect 661 1147 677 1181
rect 745 1147 761 1181
rect 661 1109 761 1147
rect 819 1181 919 1197
rect 819 1147 835 1181
rect 903 1147 919 1181
rect 819 1109 919 1147
rect -919 71 -819 109
rect -919 37 -903 71
rect -835 37 -819 71
rect -919 21 -819 37
rect -761 71 -661 109
rect -761 37 -745 71
rect -677 37 -661 71
rect -761 21 -661 37
rect -603 71 -503 109
rect -603 37 -587 71
rect -519 37 -503 71
rect -603 21 -503 37
rect -445 71 -345 109
rect -445 37 -429 71
rect -361 37 -345 71
rect -445 21 -345 37
rect -287 71 -187 109
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 109
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 109
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 109
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect 345 71 445 109
rect 345 37 361 71
rect 429 37 445 71
rect 345 21 445 37
rect 503 71 603 109
rect 503 37 519 71
rect 587 37 603 71
rect 503 21 603 37
rect 661 71 761 109
rect 661 37 677 71
rect 745 37 761 71
rect 661 21 761 37
rect 819 71 919 109
rect 819 37 835 71
rect 903 37 919 71
rect 819 21 919 37
rect -919 -37 -819 -21
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -919 -109 -819 -71
rect -761 -37 -661 -21
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -761 -109 -661 -71
rect -603 -37 -503 -21
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -603 -109 -503 -71
rect -445 -37 -345 -21
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -445 -109 -345 -71
rect -287 -37 -187 -21
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -287 -109 -187 -71
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -109 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -109 129 -71
rect 187 -37 287 -21
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 187 -109 287 -71
rect 345 -37 445 -21
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 345 -109 445 -71
rect 503 -37 603 -21
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 503 -109 603 -71
rect 661 -37 761 -21
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 661 -109 761 -71
rect 819 -37 919 -21
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 819 -109 919 -71
rect -919 -1147 -819 -1109
rect -919 -1181 -903 -1147
rect -835 -1181 -819 -1147
rect -919 -1197 -819 -1181
rect -761 -1147 -661 -1109
rect -761 -1181 -745 -1147
rect -677 -1181 -661 -1147
rect -761 -1197 -661 -1181
rect -603 -1147 -503 -1109
rect -603 -1181 -587 -1147
rect -519 -1181 -503 -1147
rect -603 -1197 -503 -1181
rect -445 -1147 -345 -1109
rect -445 -1181 -429 -1147
rect -361 -1181 -345 -1147
rect -445 -1197 -345 -1181
rect -287 -1147 -187 -1109
rect -287 -1181 -271 -1147
rect -203 -1181 -187 -1147
rect -287 -1197 -187 -1181
rect -129 -1147 -29 -1109
rect -129 -1181 -113 -1147
rect -45 -1181 -29 -1147
rect -129 -1197 -29 -1181
rect 29 -1147 129 -1109
rect 29 -1181 45 -1147
rect 113 -1181 129 -1147
rect 29 -1197 129 -1181
rect 187 -1147 287 -1109
rect 187 -1181 203 -1147
rect 271 -1181 287 -1147
rect 187 -1197 287 -1181
rect 345 -1147 445 -1109
rect 345 -1181 361 -1147
rect 429 -1181 445 -1147
rect 345 -1197 445 -1181
rect 503 -1147 603 -1109
rect 503 -1181 519 -1147
rect 587 -1181 603 -1147
rect 503 -1197 603 -1181
rect 661 -1147 761 -1109
rect 661 -1181 677 -1147
rect 745 -1181 761 -1147
rect 661 -1197 761 -1181
rect 819 -1147 919 -1109
rect 819 -1181 835 -1147
rect 903 -1181 919 -1147
rect 819 -1197 919 -1181
<< polycont >>
rect -903 1147 -835 1181
rect -745 1147 -677 1181
rect -587 1147 -519 1181
rect -429 1147 -361 1181
rect -271 1147 -203 1181
rect -113 1147 -45 1181
rect 45 1147 113 1181
rect 203 1147 271 1181
rect 361 1147 429 1181
rect 519 1147 587 1181
rect 677 1147 745 1181
rect 835 1147 903 1181
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect -903 -1181 -835 -1147
rect -745 -1181 -677 -1147
rect -587 -1181 -519 -1147
rect -429 -1181 -361 -1147
rect -271 -1181 -203 -1147
rect -113 -1181 -45 -1147
rect 45 -1181 113 -1147
rect 203 -1181 271 -1147
rect 361 -1181 429 -1147
rect 519 -1181 587 -1147
rect 677 -1181 745 -1147
rect 835 -1181 903 -1147
<< locali >>
rect -1099 1285 -1003 1319
rect 1003 1285 1099 1319
rect -1099 1223 -1065 1285
rect 1065 1223 1099 1285
rect -919 1147 -903 1181
rect -835 1147 -819 1181
rect -761 1147 -745 1181
rect -677 1147 -661 1181
rect -603 1147 -587 1181
rect -519 1147 -503 1181
rect -445 1147 -429 1181
rect -361 1147 -345 1181
rect -287 1147 -271 1181
rect -203 1147 -187 1181
rect -129 1147 -113 1181
rect -45 1147 -29 1181
rect 29 1147 45 1181
rect 113 1147 129 1181
rect 187 1147 203 1181
rect 271 1147 287 1181
rect 345 1147 361 1181
rect 429 1147 445 1181
rect 503 1147 519 1181
rect 587 1147 603 1181
rect 661 1147 677 1181
rect 745 1147 761 1181
rect 819 1147 835 1181
rect 903 1147 919 1181
rect -965 1097 -931 1113
rect -965 105 -931 121
rect -807 1097 -773 1113
rect -807 105 -773 121
rect -649 1097 -615 1113
rect -649 105 -615 121
rect -491 1097 -457 1113
rect -491 105 -457 121
rect -333 1097 -299 1113
rect -333 105 -299 121
rect -175 1097 -141 1113
rect -175 105 -141 121
rect -17 1097 17 1113
rect -17 105 17 121
rect 141 1097 175 1113
rect 141 105 175 121
rect 299 1097 333 1113
rect 299 105 333 121
rect 457 1097 491 1113
rect 457 105 491 121
rect 615 1097 649 1113
rect 615 105 649 121
rect 773 1097 807 1113
rect 773 105 807 121
rect 931 1097 965 1113
rect 931 105 965 121
rect -919 37 -903 71
rect -835 37 -819 71
rect -761 37 -745 71
rect -677 37 -661 71
rect -603 37 -587 71
rect -519 37 -503 71
rect -445 37 -429 71
rect -361 37 -345 71
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect 345 37 361 71
rect 429 37 445 71
rect 503 37 519 71
rect 587 37 603 71
rect 661 37 677 71
rect 745 37 761 71
rect 819 37 835 71
rect 903 37 919 71
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 819 -71 835 -37
rect 903 -71 919 -37
rect -965 -121 -931 -105
rect -965 -1113 -931 -1097
rect -807 -121 -773 -105
rect -807 -1113 -773 -1097
rect -649 -121 -615 -105
rect -649 -1113 -615 -1097
rect -491 -121 -457 -105
rect -491 -1113 -457 -1097
rect -333 -121 -299 -105
rect -333 -1113 -299 -1097
rect -175 -121 -141 -105
rect -175 -1113 -141 -1097
rect -17 -121 17 -105
rect -17 -1113 17 -1097
rect 141 -121 175 -105
rect 141 -1113 175 -1097
rect 299 -121 333 -105
rect 299 -1113 333 -1097
rect 457 -121 491 -105
rect 457 -1113 491 -1097
rect 615 -121 649 -105
rect 615 -1113 649 -1097
rect 773 -121 807 -105
rect 773 -1113 807 -1097
rect 931 -121 965 -105
rect 931 -1113 965 -1097
rect -919 -1181 -903 -1147
rect -835 -1181 -819 -1147
rect -761 -1181 -745 -1147
rect -677 -1181 -661 -1147
rect -603 -1181 -587 -1147
rect -519 -1181 -503 -1147
rect -445 -1181 -429 -1147
rect -361 -1181 -345 -1147
rect -287 -1181 -271 -1147
rect -203 -1181 -187 -1147
rect -129 -1181 -113 -1147
rect -45 -1181 -29 -1147
rect 29 -1181 45 -1147
rect 113 -1181 129 -1147
rect 187 -1181 203 -1147
rect 271 -1181 287 -1147
rect 345 -1181 361 -1147
rect 429 -1181 445 -1147
rect 503 -1181 519 -1147
rect 587 -1181 603 -1147
rect 661 -1181 677 -1147
rect 745 -1181 761 -1147
rect 819 -1181 835 -1147
rect 903 -1181 919 -1147
rect -1099 -1285 -1065 -1223
rect 1065 -1285 1099 -1223
rect -1099 -1319 -1003 -1285
rect 1003 -1319 1099 -1285
<< viali >>
rect -903 1147 -835 1181
rect -745 1147 -677 1181
rect -587 1147 -519 1181
rect -429 1147 -361 1181
rect -271 1147 -203 1181
rect -113 1147 -45 1181
rect 45 1147 113 1181
rect 203 1147 271 1181
rect 361 1147 429 1181
rect 519 1147 587 1181
rect 677 1147 745 1181
rect 835 1147 903 1181
rect -965 121 -931 1097
rect -807 121 -773 1097
rect -649 121 -615 1097
rect -491 121 -457 1097
rect -333 121 -299 1097
rect -175 121 -141 1097
rect -17 121 17 1097
rect 141 121 175 1097
rect 299 121 333 1097
rect 457 121 491 1097
rect 615 121 649 1097
rect 773 121 807 1097
rect 931 121 965 1097
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect -965 -1097 -931 -121
rect -807 -1097 -773 -121
rect -649 -1097 -615 -121
rect -491 -1097 -457 -121
rect -333 -1097 -299 -121
rect -175 -1097 -141 -121
rect -17 -1097 17 -121
rect 141 -1097 175 -121
rect 299 -1097 333 -121
rect 457 -1097 491 -121
rect 615 -1097 649 -121
rect 773 -1097 807 -121
rect 931 -1097 965 -121
rect -903 -1181 -835 -1147
rect -745 -1181 -677 -1147
rect -587 -1181 -519 -1147
rect -429 -1181 -361 -1147
rect -271 -1181 -203 -1147
rect -113 -1181 -45 -1147
rect 45 -1181 113 -1147
rect 203 -1181 271 -1147
rect 361 -1181 429 -1147
rect 519 -1181 587 -1147
rect 677 -1181 745 -1147
rect 835 -1181 903 -1147
<< metal1 >>
rect -915 1181 -823 1187
rect -915 1147 -903 1181
rect -835 1147 -823 1181
rect -915 1141 -823 1147
rect -757 1181 -665 1187
rect -757 1147 -745 1181
rect -677 1147 -665 1181
rect -757 1141 -665 1147
rect -599 1181 -507 1187
rect -599 1147 -587 1181
rect -519 1147 -507 1181
rect -599 1141 -507 1147
rect -441 1181 -349 1187
rect -441 1147 -429 1181
rect -361 1147 -349 1181
rect -441 1141 -349 1147
rect -283 1181 -191 1187
rect -283 1147 -271 1181
rect -203 1147 -191 1181
rect -283 1141 -191 1147
rect -125 1181 -33 1187
rect -125 1147 -113 1181
rect -45 1147 -33 1181
rect -125 1141 -33 1147
rect 33 1181 125 1187
rect 33 1147 45 1181
rect 113 1147 125 1181
rect 33 1141 125 1147
rect 191 1181 283 1187
rect 191 1147 203 1181
rect 271 1147 283 1181
rect 191 1141 283 1147
rect 349 1181 441 1187
rect 349 1147 361 1181
rect 429 1147 441 1181
rect 349 1141 441 1147
rect 507 1181 599 1187
rect 507 1147 519 1181
rect 587 1147 599 1181
rect 507 1141 599 1147
rect 665 1181 757 1187
rect 665 1147 677 1181
rect 745 1147 757 1181
rect 665 1141 757 1147
rect 823 1181 915 1187
rect 823 1147 835 1181
rect 903 1147 915 1181
rect 823 1141 915 1147
rect -971 1097 -925 1109
rect -971 121 -965 1097
rect -931 121 -925 1097
rect -971 109 -925 121
rect -813 1097 -767 1109
rect -813 121 -807 1097
rect -773 121 -767 1097
rect -813 109 -767 121
rect -655 1097 -609 1109
rect -655 121 -649 1097
rect -615 121 -609 1097
rect -655 109 -609 121
rect -497 1097 -451 1109
rect -497 121 -491 1097
rect -457 121 -451 1097
rect -497 109 -451 121
rect -339 1097 -293 1109
rect -339 121 -333 1097
rect -299 121 -293 1097
rect -339 109 -293 121
rect -181 1097 -135 1109
rect -181 121 -175 1097
rect -141 121 -135 1097
rect -181 109 -135 121
rect -23 1097 23 1109
rect -23 121 -17 1097
rect 17 121 23 1097
rect -23 109 23 121
rect 135 1097 181 1109
rect 135 121 141 1097
rect 175 121 181 1097
rect 135 109 181 121
rect 293 1097 339 1109
rect 293 121 299 1097
rect 333 121 339 1097
rect 293 109 339 121
rect 451 1097 497 1109
rect 451 121 457 1097
rect 491 121 497 1097
rect 451 109 497 121
rect 609 1097 655 1109
rect 609 121 615 1097
rect 649 121 655 1097
rect 609 109 655 121
rect 767 1097 813 1109
rect 767 121 773 1097
rect 807 121 813 1097
rect 767 109 813 121
rect 925 1097 971 1109
rect 925 121 931 1097
rect 965 121 971 1097
rect 925 109 971 121
rect -915 71 -823 77
rect -915 37 -903 71
rect -835 37 -823 71
rect -915 31 -823 37
rect -757 71 -665 77
rect -757 37 -745 71
rect -677 37 -665 71
rect -757 31 -665 37
rect -599 71 -507 77
rect -599 37 -587 71
rect -519 37 -507 71
rect -599 31 -507 37
rect -441 71 -349 77
rect -441 37 -429 71
rect -361 37 -349 71
rect -441 31 -349 37
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect 349 71 441 77
rect 349 37 361 71
rect 429 37 441 71
rect 349 31 441 37
rect 507 71 599 77
rect 507 37 519 71
rect 587 37 599 71
rect 507 31 599 37
rect 665 71 757 77
rect 665 37 677 71
rect 745 37 757 71
rect 665 31 757 37
rect 823 71 915 77
rect 823 37 835 71
rect 903 37 915 71
rect 823 31 915 37
rect -915 -37 -823 -31
rect -915 -71 -903 -37
rect -835 -71 -823 -37
rect -915 -77 -823 -71
rect -757 -37 -665 -31
rect -757 -71 -745 -37
rect -677 -71 -665 -37
rect -757 -77 -665 -71
rect -599 -37 -507 -31
rect -599 -71 -587 -37
rect -519 -71 -507 -37
rect -599 -77 -507 -71
rect -441 -37 -349 -31
rect -441 -71 -429 -37
rect -361 -71 -349 -37
rect -441 -77 -349 -71
rect -283 -37 -191 -31
rect -283 -71 -271 -37
rect -203 -71 -191 -37
rect -283 -77 -191 -71
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect 191 -37 283 -31
rect 191 -71 203 -37
rect 271 -71 283 -37
rect 191 -77 283 -71
rect 349 -37 441 -31
rect 349 -71 361 -37
rect 429 -71 441 -37
rect 349 -77 441 -71
rect 507 -37 599 -31
rect 507 -71 519 -37
rect 587 -71 599 -37
rect 507 -77 599 -71
rect 665 -37 757 -31
rect 665 -71 677 -37
rect 745 -71 757 -37
rect 665 -77 757 -71
rect 823 -37 915 -31
rect 823 -71 835 -37
rect 903 -71 915 -37
rect 823 -77 915 -71
rect -971 -121 -925 -109
rect -971 -1097 -965 -121
rect -931 -1097 -925 -121
rect -971 -1109 -925 -1097
rect -813 -121 -767 -109
rect -813 -1097 -807 -121
rect -773 -1097 -767 -121
rect -813 -1109 -767 -1097
rect -655 -121 -609 -109
rect -655 -1097 -649 -121
rect -615 -1097 -609 -121
rect -655 -1109 -609 -1097
rect -497 -121 -451 -109
rect -497 -1097 -491 -121
rect -457 -1097 -451 -121
rect -497 -1109 -451 -1097
rect -339 -121 -293 -109
rect -339 -1097 -333 -121
rect -299 -1097 -293 -121
rect -339 -1109 -293 -1097
rect -181 -121 -135 -109
rect -181 -1097 -175 -121
rect -141 -1097 -135 -121
rect -181 -1109 -135 -1097
rect -23 -121 23 -109
rect -23 -1097 -17 -121
rect 17 -1097 23 -121
rect -23 -1109 23 -1097
rect 135 -121 181 -109
rect 135 -1097 141 -121
rect 175 -1097 181 -121
rect 135 -1109 181 -1097
rect 293 -121 339 -109
rect 293 -1097 299 -121
rect 333 -1097 339 -121
rect 293 -1109 339 -1097
rect 451 -121 497 -109
rect 451 -1097 457 -121
rect 491 -1097 497 -121
rect 451 -1109 497 -1097
rect 609 -121 655 -109
rect 609 -1097 615 -121
rect 649 -1097 655 -121
rect 609 -1109 655 -1097
rect 767 -121 813 -109
rect 767 -1097 773 -121
rect 807 -1097 813 -121
rect 767 -1109 813 -1097
rect 925 -121 971 -109
rect 925 -1097 931 -121
rect 965 -1097 971 -121
rect 925 -1109 971 -1097
rect -915 -1147 -823 -1141
rect -915 -1181 -903 -1147
rect -835 -1181 -823 -1147
rect -915 -1187 -823 -1181
rect -757 -1147 -665 -1141
rect -757 -1181 -745 -1147
rect -677 -1181 -665 -1147
rect -757 -1187 -665 -1181
rect -599 -1147 -507 -1141
rect -599 -1181 -587 -1147
rect -519 -1181 -507 -1147
rect -599 -1187 -507 -1181
rect -441 -1147 -349 -1141
rect -441 -1181 -429 -1147
rect -361 -1181 -349 -1147
rect -441 -1187 -349 -1181
rect -283 -1147 -191 -1141
rect -283 -1181 -271 -1147
rect -203 -1181 -191 -1147
rect -283 -1187 -191 -1181
rect -125 -1147 -33 -1141
rect -125 -1181 -113 -1147
rect -45 -1181 -33 -1147
rect -125 -1187 -33 -1181
rect 33 -1147 125 -1141
rect 33 -1181 45 -1147
rect 113 -1181 125 -1147
rect 33 -1187 125 -1181
rect 191 -1147 283 -1141
rect 191 -1181 203 -1147
rect 271 -1181 283 -1147
rect 191 -1187 283 -1181
rect 349 -1147 441 -1141
rect 349 -1181 361 -1147
rect 429 -1181 441 -1147
rect 349 -1187 441 -1181
rect 507 -1147 599 -1141
rect 507 -1181 519 -1147
rect 587 -1181 599 -1147
rect 507 -1187 599 -1181
rect 665 -1147 757 -1141
rect 665 -1181 677 -1147
rect 745 -1181 757 -1147
rect 665 -1187 757 -1181
rect 823 -1147 915 -1141
rect 823 -1181 835 -1147
rect 903 -1181 915 -1147
rect 823 -1187 915 -1181
<< properties >>
string FIXED_BBOX -1082 -1302 1082 1302
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.50 m 2 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
