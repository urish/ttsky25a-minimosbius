magic
tech sky130A
magscale 1 2
timestamp 1757283573
<< nwell >>
rect -146 7546 390 7868
rect 252 6704 258 6778
rect 252 5616 258 5690
rect 1832 4766 1900 4849
rect 252 4528 258 4602
<< pwell >>
rect 1865 4907 1900 4912
<< pdiff >>
rect 1852 4766 1900 4813
<< locali >>
rect 1841 4894 1891 4912
rect 1841 4788 1848 4894
rect 1882 4788 1891 4894
rect 1841 4766 1891 4788
<< viali >>
rect 96 7368 130 7546
rect 228 7438 334 7544
rect 3318 7104 3352 7138
rect 1754 6970 1788 7004
rect 3594 6970 3628 7004
rect 10 6830 44 6936
rect 1500 6828 1534 6862
rect 1852 6828 1886 6862
rect 1764 6622 1798 6656
rect 2116 6622 2150 6656
rect 20 6480 54 6514
rect 1860 6480 1894 6514
rect 3604 6502 3638 6608
rect 298 6332 332 6366
rect 3318 6026 3352 6060
rect 1754 5882 1788 5916
rect 3594 5882 3628 5916
rect 10 5742 44 5848
rect 1500 5740 1534 5774
rect 1852 5740 1886 5774
rect 1764 5534 1798 5568
rect 20 5392 54 5426
rect 298 5244 332 5278
rect 1764 5234 1798 5268
rect 8 4788 42 4894
rect 182 4852 216 4886
rect 296 4854 330 4888
rect 468 4788 502 4894
rect 642 4852 676 4886
rect 756 4854 790 4888
rect 928 4788 962 4894
rect 1102 4852 1136 4886
rect 1216 4854 1250 4888
rect 1388 4788 1422 4894
rect 1562 4852 1596 4886
rect 1676 4854 1710 4888
rect 1848 4788 1882 4894
rect 2022 4852 2056 4886
rect 2136 4854 2170 4888
rect 2308 4788 2342 4894
rect 2482 4852 2516 4886
rect 2596 4854 2630 4888
rect 2768 4788 2802 4894
rect 2942 4852 2976 4886
rect 3056 4854 3090 4888
<< metal1 >>
rect -102 7854 232 7858
rect -102 7802 50 7854
rect 230 7802 236 7854
rect -102 7788 232 7802
rect 18 7548 146 7556
rect 18 7432 24 7548
rect 140 7432 146 7548
rect 18 7426 96 7432
rect 84 7368 96 7426
rect 130 7426 146 7432
rect 216 7544 346 7554
rect 216 7438 228 7544
rect 334 7500 346 7544
rect 1040 7508 1168 7514
rect 1040 7500 1046 7508
rect 334 7460 1046 7500
rect 334 7438 346 7460
rect 1040 7456 1046 7460
rect 1162 7500 1168 7508
rect 1802 7506 1930 7512
rect 1802 7500 1808 7506
rect 1162 7460 1808 7500
rect 1162 7456 1168 7460
rect 1040 7450 1168 7456
rect 1802 7454 1808 7460
rect 1924 7500 1930 7506
rect 3502 7506 3630 7512
rect 3502 7500 3508 7506
rect 1924 7460 3508 7500
rect 1924 7454 1930 7460
rect 1802 7448 1930 7454
rect 3502 7454 3508 7460
rect 3624 7454 3630 7506
rect 3502 7448 3630 7454
rect 216 7426 346 7438
rect 130 7368 142 7426
rect 84 7362 142 7368
rect 802 7424 930 7430
rect 802 7372 808 7424
rect 924 7418 930 7424
rect 2578 7424 2706 7430
rect 2578 7418 2584 7424
rect 924 7378 2584 7418
rect 924 7372 930 7378
rect 802 7366 930 7372
rect 2578 7372 2584 7378
rect 2700 7372 2706 7424
rect 2578 7366 2706 7372
rect 364 7258 370 7310
rect 550 7258 556 7310
rect 802 7160 866 7166
rect 802 7108 808 7160
rect 860 7108 866 7160
rect 802 7102 866 7108
rect 2642 7160 2706 7166
rect 2642 7108 2648 7160
rect 2700 7108 2706 7160
rect 2642 7102 2706 7108
rect 3302 7154 3368 7160
rect 3302 7100 3308 7154
rect 3362 7100 3368 7154
rect 3302 7094 3368 7100
rect 1738 7004 1802 7010
rect 1738 6952 1744 7004
rect 1796 6952 1802 7004
rect 4 6936 50 6948
rect 1738 6946 1802 6952
rect 3578 7004 3642 7010
rect 3578 6952 3584 7004
rect 3636 6952 3642 7004
rect 3578 6946 3642 6952
rect 4 6830 10 6936
rect 44 6890 50 6936
rect 282 6898 346 6904
rect 282 6890 288 6898
rect 44 6854 288 6890
rect 44 6830 50 6854
rect 282 6846 288 6854
rect 340 6846 346 6898
rect 1680 6878 1744 6884
rect 282 6840 346 6846
rect 1488 6862 1552 6868
rect 4 6818 50 6830
rect 1488 6828 1500 6862
rect 1534 6860 1552 6862
rect 1680 6860 1686 6878
rect 1534 6830 1686 6860
rect 1534 6828 1552 6830
rect 1488 6822 1552 6828
rect 1680 6826 1686 6830
rect 1738 6860 1744 6878
rect 1840 6862 1898 6868
rect 1840 6860 1852 6862
rect 1738 6830 1852 6860
rect 1738 6826 1744 6830
rect 1680 6820 1744 6826
rect 1840 6828 1852 6830
rect 1886 6828 1898 6862
rect 1840 6822 1898 6828
rect 44 6714 50 6766
rect 230 6714 236 6766
rect 1648 6656 1712 6662
rect 1648 6604 1654 6656
rect 1706 6654 1712 6656
rect 1752 6656 1810 6662
rect 1752 6654 1764 6656
rect 1706 6624 1764 6654
rect 1706 6604 1712 6624
rect 1752 6622 1764 6624
rect 1798 6654 1810 6656
rect 2098 6656 2162 6662
rect 2098 6654 2116 6656
rect 1798 6624 2116 6654
rect 1798 6622 1810 6624
rect 1752 6616 1810 6622
rect 2098 6622 2116 6624
rect 2150 6622 2162 6656
rect 2098 6616 2162 6622
rect 1648 6598 1712 6604
rect 3598 6608 3644 6620
rect 3302 6582 3366 6588
rect 4 6532 68 6538
rect 4 6480 10 6532
rect 62 6480 68 6532
rect 4 6474 68 6480
rect 1844 6532 1908 6538
rect 1844 6480 1850 6532
rect 1902 6480 1908 6532
rect 3302 6530 3308 6582
rect 3360 6576 3366 6582
rect 3598 6576 3604 6608
rect 3360 6536 3604 6576
rect 3360 6530 3366 6536
rect 3302 6524 3366 6530
rect 3598 6502 3604 6536
rect 3638 6502 3644 6608
rect 3598 6490 3644 6502
rect 1844 6474 1908 6480
rect 804 6386 868 6392
rect 282 6374 346 6380
rect 282 6322 288 6374
rect 340 6322 346 6374
rect 804 6334 810 6386
rect 862 6334 868 6386
rect 804 6328 868 6334
rect 2644 6386 2708 6392
rect 2644 6334 2650 6386
rect 2702 6334 2708 6386
rect 2644 6328 2708 6334
rect 282 6316 346 6322
rect 364 6170 370 6222
rect 550 6170 556 6222
rect 802 6072 866 6078
rect 802 6020 808 6072
rect 860 6020 866 6072
rect 802 6014 866 6020
rect 2642 6072 2706 6078
rect 2642 6020 2648 6072
rect 2700 6020 2706 6072
rect 2642 6014 2706 6020
rect 3302 6068 3366 6074
rect 3302 6016 3308 6068
rect 3360 6016 3366 6068
rect 3302 6010 3366 6016
rect 1738 5916 1802 5922
rect 1738 5864 1744 5916
rect 1796 5864 1802 5916
rect 4 5848 50 5860
rect 1738 5858 1802 5864
rect 3578 5916 3642 5922
rect 3578 5864 3584 5916
rect 3636 5864 3642 5916
rect 3578 5858 3642 5864
rect 4 5742 10 5848
rect 44 5802 50 5848
rect 282 5810 346 5816
rect 282 5802 288 5810
rect 44 5766 288 5802
rect 44 5742 50 5766
rect 282 5758 288 5766
rect 340 5758 346 5810
rect 2120 5794 2184 5800
rect 282 5752 346 5758
rect 1488 5774 1552 5780
rect 4 5730 50 5742
rect 1488 5740 1500 5774
rect 1534 5772 1552 5774
rect 1840 5774 1898 5780
rect 1840 5772 1852 5774
rect 1534 5742 1852 5772
rect 1534 5740 1552 5742
rect 1488 5734 1552 5740
rect 1840 5740 1852 5742
rect 1886 5772 1898 5774
rect 2120 5772 2126 5794
rect 1886 5742 2126 5772
rect 2178 5742 2184 5794
rect 1886 5740 1898 5742
rect 1840 5734 1898 5740
rect 2120 5736 2184 5742
rect 44 5626 70 5678
rect 230 5626 236 5678
rect 1752 5568 1810 5574
rect 1752 5534 1764 5568
rect 1798 5534 1810 5568
rect 4 5444 68 5450
rect 4 5392 10 5444
rect 62 5392 68 5444
rect 4 5386 68 5392
rect 802 5298 866 5304
rect 282 5286 346 5292
rect 282 5234 288 5286
rect 340 5234 346 5286
rect 802 5246 808 5298
rect 862 5246 866 5298
rect 802 5240 866 5246
rect 1752 5268 1810 5534
rect 3406 5292 3534 5298
rect 2460 5276 2524 5282
rect 2460 5268 2466 5276
rect 282 5228 346 5234
rect 1752 5234 1764 5268
rect 1798 5234 2466 5268
rect 1752 5228 1810 5234
rect 2460 5224 2466 5234
rect 2518 5268 2524 5276
rect 3406 5268 3412 5292
rect 2518 5240 3412 5268
rect 3528 5240 3534 5292
rect 2518 5234 3534 5240
rect 2518 5224 2524 5234
rect 2460 5218 2524 5224
rect 364 5082 370 5134
rect 550 5082 556 5134
rect 3186 5062 3702 5158
rect 2258 5020 2386 5026
rect 2258 5014 2264 5020
rect 2018 5012 2264 5014
rect 642 5006 706 5012
rect 642 4954 648 5006
rect 700 5000 706 5006
rect 700 4960 794 5000
rect 700 4954 706 4960
rect 642 4948 706 4954
rect -6 4898 58 4904
rect -6 4782 0 4898
rect 52 4782 58 4898
rect -6 4776 58 4782
rect 176 4886 222 4898
rect 176 4852 182 4886
rect 216 4852 222 4886
rect 176 4716 222 4852
rect 282 4896 346 4902
rect 282 4844 288 4896
rect 340 4844 346 4896
rect 282 4838 346 4844
rect 454 4898 518 4904
rect 754 4902 794 4960
rect 2016 4974 2264 5012
rect 454 4782 460 4898
rect 512 4782 518 4898
rect 454 4776 518 4782
rect 636 4886 682 4898
rect 636 4852 642 4886
rect 676 4852 682 4886
rect 636 4716 682 4852
rect 742 4896 806 4902
rect 742 4844 748 4896
rect 800 4844 806 4896
rect 742 4838 806 4844
rect 914 4898 978 4904
rect 914 4782 920 4898
rect 972 4782 978 4898
rect 914 4776 978 4782
rect 1096 4886 1142 4898
rect 1096 4852 1102 4886
rect 1136 4852 1142 4886
rect 1096 4716 1142 4852
rect 1202 4896 1266 4902
rect 1202 4844 1208 4896
rect 1260 4844 1266 4896
rect 1202 4838 1266 4844
rect 1374 4898 1438 4904
rect 1374 4782 1380 4898
rect 1432 4782 1438 4898
rect 1374 4776 1438 4782
rect 1556 4886 1602 4898
rect 1556 4852 1562 4886
rect 1596 4852 1602 4886
rect 1556 4716 1602 4852
rect 1662 4896 1726 4902
rect 1662 4844 1668 4896
rect 1720 4844 1726 4896
rect 1662 4838 1726 4844
rect 1834 4898 1898 4904
rect 1834 4782 1840 4898
rect 1892 4782 1898 4898
rect 1834 4776 1898 4782
rect 2016 4886 2062 4974
rect 2258 4968 2264 4974
rect 2380 5014 2386 5020
rect 2380 4974 2522 5014
rect 2380 4968 2386 4974
rect 2258 4962 2386 4968
rect 2016 4852 2022 4886
rect 2056 4852 2062 4886
rect 2016 4716 2062 4852
rect 2122 4896 2186 4902
rect 2122 4844 2128 4896
rect 2180 4844 2186 4896
rect 2122 4838 2186 4844
rect 2294 4898 2358 4904
rect 2294 4782 2300 4898
rect 2352 4782 2358 4898
rect 2294 4776 2358 4782
rect 2476 4886 2522 4974
rect 2476 4852 2482 4886
rect 2516 4852 2522 4886
rect 2476 4716 2522 4852
rect 2582 4896 2646 4902
rect 2582 4844 2588 4896
rect 2640 4844 2646 4896
rect 2582 4838 2646 4844
rect 2754 4898 2818 4904
rect 2754 4782 2760 4898
rect 2812 4782 2818 4898
rect 2754 4776 2818 4782
rect 2936 4886 2982 4898
rect 2936 4852 2942 4886
rect 2976 4852 2982 4886
rect 2936 4716 2982 4852
rect 3042 4896 3106 4902
rect 3042 4844 3048 4896
rect 3100 4844 3106 4896
rect 3042 4838 3106 4844
rect -66 4676 3716 4716
rect 44 4538 50 4590
rect 230 4538 236 4590
rect 3198 4518 3714 4614
rect 2066 -23168 2130 -23162
rect 2066 -23196 2072 -23168
rect 890 -23256 2072 -23196
rect 890 -23436 950 -23256
rect 2066 -23284 2072 -23256
rect 2124 -23196 2130 -23168
rect 2124 -23256 2132 -23196
rect 2124 -23284 2130 -23256
rect 2066 -23290 2130 -23284
<< via1 >>
rect 50 7802 230 7854
rect 24 7546 140 7548
rect 24 7432 96 7546
rect 96 7432 130 7546
rect 130 7432 140 7546
rect 1046 7456 1162 7508
rect 1808 7454 1924 7506
rect 3508 7454 3624 7506
rect 808 7372 924 7424
rect 2584 7372 2700 7424
rect 370 7258 550 7310
rect 808 7108 860 7160
rect 2648 7108 2700 7160
rect 3308 7138 3362 7154
rect 3308 7104 3318 7138
rect 3318 7104 3352 7138
rect 3352 7104 3362 7138
rect 3308 7100 3362 7104
rect 1744 6970 1754 7004
rect 1754 6970 1788 7004
rect 1788 6970 1796 7004
rect 1744 6952 1796 6970
rect 3584 6970 3594 7004
rect 3594 6970 3628 7004
rect 3628 6970 3636 7004
rect 3584 6952 3636 6970
rect 288 6846 340 6898
rect 1686 6826 1738 6878
rect 50 6714 230 6766
rect 1654 6604 1706 6656
rect 10 6514 62 6532
rect 10 6480 20 6514
rect 20 6480 54 6514
rect 54 6480 62 6514
rect 1850 6514 1902 6532
rect 1850 6480 1860 6514
rect 1860 6480 1894 6514
rect 1894 6480 1902 6514
rect 3308 6530 3360 6582
rect 288 6366 340 6374
rect 288 6332 298 6366
rect 298 6332 332 6366
rect 332 6332 340 6366
rect 288 6322 340 6332
rect 810 6334 862 6386
rect 2650 6334 2702 6386
rect 370 6170 550 6222
rect 808 6020 860 6072
rect 2648 6020 2700 6072
rect 3308 6060 3360 6068
rect 3308 6026 3318 6060
rect 3318 6026 3352 6060
rect 3352 6026 3360 6060
rect 3308 6016 3360 6026
rect 1744 5882 1754 5916
rect 1754 5882 1788 5916
rect 1788 5882 1796 5916
rect 1744 5864 1796 5882
rect 3584 5882 3594 5916
rect 3594 5882 3628 5916
rect 3628 5882 3636 5916
rect 3584 5864 3636 5882
rect 288 5758 340 5810
rect 2126 5742 2178 5794
rect 70 5626 230 5678
rect 10 5426 62 5444
rect 10 5392 20 5426
rect 20 5392 54 5426
rect 54 5392 62 5426
rect 288 5278 340 5286
rect 288 5244 298 5278
rect 298 5244 332 5278
rect 332 5244 340 5278
rect 288 5234 340 5244
rect 808 5246 862 5298
rect 2466 5224 2518 5276
rect 3412 5240 3528 5292
rect 370 5082 550 5134
rect 648 4954 700 5006
rect 0 4894 52 4898
rect 0 4788 8 4894
rect 8 4788 42 4894
rect 42 4788 52 4894
rect 0 4782 52 4788
rect 288 4888 340 4896
rect 288 4854 296 4888
rect 296 4854 330 4888
rect 330 4854 340 4888
rect 288 4844 340 4854
rect 460 4894 512 4898
rect 460 4788 468 4894
rect 468 4788 502 4894
rect 502 4788 512 4894
rect 460 4782 512 4788
rect 748 4888 800 4896
rect 748 4854 756 4888
rect 756 4854 790 4888
rect 790 4854 800 4888
rect 748 4844 800 4854
rect 920 4894 972 4898
rect 920 4788 928 4894
rect 928 4788 962 4894
rect 962 4788 972 4894
rect 920 4782 972 4788
rect 1208 4888 1260 4896
rect 1208 4854 1216 4888
rect 1216 4854 1250 4888
rect 1250 4854 1260 4888
rect 1208 4844 1260 4854
rect 1380 4894 1432 4898
rect 1380 4788 1388 4894
rect 1388 4788 1422 4894
rect 1422 4788 1432 4894
rect 1380 4782 1432 4788
rect 1668 4888 1720 4896
rect 1668 4854 1676 4888
rect 1676 4854 1710 4888
rect 1710 4854 1720 4888
rect 1668 4844 1720 4854
rect 1840 4894 1892 4898
rect 1840 4788 1848 4894
rect 1848 4788 1882 4894
rect 1882 4788 1892 4894
rect 1840 4782 1892 4788
rect 2264 4968 2380 5020
rect 2128 4888 2180 4896
rect 2128 4854 2136 4888
rect 2136 4854 2170 4888
rect 2170 4854 2180 4888
rect 2128 4844 2180 4854
rect 2300 4894 2352 4898
rect 2300 4788 2308 4894
rect 2308 4788 2342 4894
rect 2342 4788 2352 4894
rect 2300 4782 2352 4788
rect 2588 4888 2640 4896
rect 2588 4854 2596 4888
rect 2596 4854 2630 4888
rect 2630 4854 2640 4888
rect 2588 4844 2640 4854
rect 2760 4894 2812 4898
rect 2760 4788 2768 4894
rect 2768 4788 2802 4894
rect 2802 4788 2812 4894
rect 2760 4782 2812 4788
rect 3048 4888 3100 4896
rect 3048 4854 3056 4888
rect 3056 4854 3090 4888
rect 3090 4854 3100 4888
rect 3048 4844 3100 4854
rect 50 4538 230 4590
rect 2072 -23284 2124 -23168
<< metal2 >>
rect 2246 7958 2256 8014
rect 2392 7958 2402 8014
rect 22 7800 32 7856
rect 248 7800 258 7856
rect 766 7674 902 7684
rect 766 7608 902 7618
rect 14 7548 150 7558
rect 814 7430 854 7608
rect 1040 7508 1168 7514
rect 1040 7456 1046 7508
rect 1162 7456 1168 7508
rect 1040 7450 1168 7456
rect 1802 7506 1930 7512
rect 1802 7454 1808 7506
rect 1924 7454 1930 7506
rect 14 7402 150 7412
rect 802 7424 930 7430
rect 802 7372 808 7424
rect 924 7372 930 7424
rect 802 7366 930 7372
rect 342 7256 352 7312
rect 568 7256 578 7312
rect 814 7166 854 7366
rect 802 7160 866 7166
rect 802 7108 808 7160
rect 860 7108 866 7160
rect 802 7102 866 7108
rect 282 6898 346 6904
rect 282 6846 288 6898
rect 340 6846 346 6898
rect 282 6840 346 6846
rect 22 6712 32 6768
rect 248 6712 258 6768
rect 4 6534 68 6544
rect 4 6478 8 6534
rect 64 6478 68 6534
rect 4 6468 68 6478
rect 294 6380 334 6840
rect 814 6392 854 7102
rect 1088 6544 1128 7450
rect 1802 7448 1930 7454
rect 1802 7010 1842 7448
rect 1738 7004 1842 7010
rect 1738 6952 1744 7004
rect 1796 6952 1842 7004
rect 1738 6946 1842 6952
rect 1680 6878 1744 6884
rect 1680 6872 1686 6878
rect 1214 6832 1686 6872
rect 1076 6534 1140 6544
rect 1076 6478 1080 6534
rect 1136 6478 1140 6534
rect 1076 6468 1140 6478
rect 804 6386 868 6392
rect 282 6374 346 6380
rect 282 6322 288 6374
rect 340 6368 346 6374
rect 340 6328 694 6368
rect 804 6334 810 6386
rect 862 6334 868 6386
rect 804 6328 868 6334
rect 340 6322 346 6328
rect 282 6316 346 6322
rect 342 6168 352 6224
rect 568 6168 578 6224
rect 282 5810 346 5816
rect 282 5758 288 5810
rect 340 5758 346 5810
rect 282 5752 346 5758
rect 60 5624 70 5680
rect 248 5624 258 5680
rect 4 5446 68 5456
rect 4 5390 8 5446
rect 64 5390 68 5446
rect 4 5380 68 5390
rect 294 5292 334 5752
rect 282 5286 346 5292
rect 282 5280 288 5286
rect 214 5240 288 5280
rect 214 5012 254 5240
rect 282 5234 288 5240
rect 340 5234 346 5286
rect 282 5228 346 5234
rect 342 5080 352 5136
rect 568 5080 578 5136
rect 654 5012 694 6328
rect 814 6078 854 6328
rect 802 6072 866 6078
rect 802 6020 808 6072
rect 860 6020 866 6072
rect 802 6014 866 6020
rect 814 5304 854 6014
rect 1088 5452 1128 6468
rect 1074 5442 1138 5452
rect 1074 5386 1078 5442
rect 1134 5386 1138 5442
rect 1074 5376 1138 5386
rect 802 5298 866 5304
rect 802 5246 808 5298
rect 862 5246 866 5298
rect 802 5240 866 5246
rect 214 4972 334 5012
rect -6 4906 58 4916
rect -6 4772 -2 4906
rect 54 4772 58 4906
rect 294 4902 334 4972
rect 642 5006 706 5012
rect 642 4954 648 5006
rect 700 4954 706 5006
rect 642 4948 706 4954
rect 454 4906 518 4916
rect 282 4896 346 4902
rect 282 4844 288 4896
rect 340 4844 346 4896
rect 282 4838 346 4844
rect -6 4762 58 4772
rect 454 4772 458 4906
rect 514 4772 518 4906
rect 742 4896 806 4902
rect 742 4844 748 4896
rect 800 4844 806 4896
rect 742 4838 806 4844
rect 914 4898 978 4904
rect 1214 4902 1254 6832
rect 1680 6826 1686 6832
rect 1738 6826 1744 6878
rect 1680 6820 1744 6826
rect 1648 6656 1712 6662
rect 1648 6604 1654 6656
rect 1706 6604 1712 6656
rect 1648 6598 1712 6604
rect 914 4782 920 4898
rect 972 4782 978 4898
rect 1202 4896 1266 4902
rect 1202 4844 1208 4896
rect 1260 4844 1266 4896
rect 1202 4838 1266 4844
rect 1374 4898 1438 4904
rect 914 4776 978 4782
rect 1374 4782 1380 4898
rect 1432 4782 1438 4898
rect 1662 4902 1702 6598
rect 1802 6538 1842 6946
rect 1802 6532 1908 6538
rect 1802 6480 1850 6532
rect 1902 6480 1908 6532
rect 1802 6474 1908 6480
rect 1802 5922 1842 6474
rect 1738 5916 1842 5922
rect 1738 5864 1744 5916
rect 1796 5864 1842 5916
rect 1738 5858 1842 5864
rect 2120 5794 2184 5800
rect 2120 5742 2126 5794
rect 2178 5742 2184 5794
rect 2120 5736 2184 5742
rect 1828 4906 1904 4912
rect 1662 4896 1726 4902
rect 1662 4844 1668 4896
rect 1720 4844 1726 4896
rect 1662 4838 1726 4844
rect 1374 4776 1438 4782
rect 454 4762 518 4772
rect 22 4536 32 4592
rect 248 4536 258 4592
rect 926 4286 966 4776
rect 1180 4652 1220 4658
rect 1386 4652 1426 4776
rect 1828 4772 1838 4906
rect 1894 4772 1904 4906
rect 2134 4902 2174 5736
rect 2304 5026 2344 7958
rect 3502 7506 3630 7512
rect 3502 7454 3508 7506
rect 3624 7454 3630 7506
rect 3502 7448 3630 7454
rect 2578 7424 2706 7430
rect 2578 7372 2584 7424
rect 2700 7372 2706 7424
rect 2578 7366 2706 7372
rect 2654 7166 2694 7366
rect 2642 7160 2706 7166
rect 2642 7108 2648 7160
rect 2700 7108 2706 7160
rect 3302 7156 3368 7160
rect 3452 7156 3492 7160
rect 2642 7102 2706 7108
rect 2654 6392 2694 7102
rect 3296 7100 3306 7156
rect 3362 7100 3372 7156
rect 3434 7100 3444 7156
rect 3500 7100 3510 7156
rect 3302 7094 3368 7100
rect 3302 6582 3366 6588
rect 3302 6530 3308 6582
rect 3360 6530 3366 6582
rect 3302 6524 3366 6530
rect 2644 6386 2708 6392
rect 2644 6334 2650 6386
rect 2702 6334 2708 6386
rect 2644 6328 2708 6334
rect 2654 6078 2694 6328
rect 2642 6072 2706 6078
rect 3314 6074 3354 6524
rect 2642 6020 2648 6072
rect 2700 6020 2706 6072
rect 3302 6068 3366 6074
rect 3302 6062 3308 6068
rect 2642 6014 2706 6020
rect 3054 6022 3308 6062
rect 2460 5276 2524 5282
rect 2460 5224 2466 5276
rect 2518 5224 2524 5276
rect 2460 5218 2524 5224
rect 2258 5020 2386 5026
rect 2258 4968 2264 5020
rect 2380 4968 2386 5020
rect 2258 4962 2386 4968
rect 2122 4896 2186 4902
rect 2122 4844 2128 4896
rect 2180 4844 2186 4896
rect 2122 4838 2186 4844
rect 2294 4898 2358 4904
rect 2294 4782 2300 4898
rect 2352 4782 2358 4898
rect 2472 4890 2512 5218
rect 2582 4896 2646 4902
rect 2582 4890 2588 4896
rect 2472 4850 2588 4890
rect 2582 4844 2588 4850
rect 2640 4844 2646 4896
rect 2582 4838 2646 4844
rect 2754 4898 2818 4904
rect 3054 4902 3094 6022
rect 3302 6016 3308 6022
rect 3360 6016 3366 6068
rect 3302 6010 3366 6016
rect 3452 5298 3492 7100
rect 3590 7010 3630 7448
rect 3578 7004 3642 7010
rect 3578 6952 3584 7004
rect 3636 6952 3642 7004
rect 3578 6946 3642 6952
rect 3590 5922 3630 6946
rect 3578 5916 3642 5922
rect 3578 5864 3584 5916
rect 3636 5864 3642 5916
rect 3578 5858 3642 5864
rect 3406 5292 3534 5298
rect 3406 5240 3412 5292
rect 3528 5240 3534 5292
rect 3406 5234 3534 5240
rect 2294 4776 2358 4782
rect 2754 4782 2760 4898
rect 2812 4782 2818 4898
rect 3042 4896 3106 4902
rect 3042 4844 3048 4896
rect 3100 4844 3106 4896
rect 3042 4838 3106 4844
rect 2754 4776 2818 4782
rect 1828 4766 1904 4772
rect 1160 4518 1170 4652
rect 1226 4612 1426 4652
rect 1226 4518 1236 4612
rect 1180 4458 1220 4518
rect 2070 4474 2126 4484
rect 2306 4428 2346 4776
rect 2766 4654 2806 4776
rect 2758 4644 2814 4654
rect 2758 4500 2814 4510
rect 2126 4388 2346 4428
rect 2070 4328 2126 4338
rect 2060 -23294 2070 -23158
rect 2126 -23294 2136 -23158
<< via2 >>
rect 2256 7958 2392 8014
rect 32 7854 248 7856
rect 32 7802 50 7854
rect 50 7802 230 7854
rect 230 7802 248 7854
rect 32 7800 248 7802
rect 766 7618 902 7674
rect 14 7432 24 7548
rect 24 7432 140 7548
rect 140 7432 150 7548
rect 14 7412 150 7432
rect 352 7310 568 7312
rect 352 7258 370 7310
rect 370 7258 550 7310
rect 550 7258 568 7310
rect 352 7256 568 7258
rect 32 6766 248 6768
rect 32 6714 50 6766
rect 50 6714 230 6766
rect 230 6714 248 6766
rect 32 6712 248 6714
rect 8 6532 64 6534
rect 8 6480 10 6532
rect 10 6480 62 6532
rect 62 6480 64 6532
rect 8 6478 64 6480
rect 1080 6478 1136 6534
rect 352 6222 568 6224
rect 352 6170 370 6222
rect 370 6170 550 6222
rect 550 6170 568 6222
rect 352 6168 568 6170
rect 70 5678 248 5680
rect 70 5626 230 5678
rect 230 5626 248 5678
rect 70 5624 248 5626
rect 8 5444 64 5446
rect 8 5392 10 5444
rect 10 5392 62 5444
rect 62 5392 64 5444
rect 8 5390 64 5392
rect 352 5134 568 5136
rect 352 5082 370 5134
rect 370 5082 550 5134
rect 550 5082 568 5134
rect 352 5080 568 5082
rect 1078 5386 1134 5442
rect -2 4898 54 4906
rect -2 4782 0 4898
rect 0 4782 52 4898
rect 52 4782 54 4898
rect -2 4772 54 4782
rect 458 4898 514 4906
rect 458 4782 460 4898
rect 460 4782 512 4898
rect 512 4782 514 4898
rect 458 4772 514 4782
rect 32 4590 248 4592
rect 32 4538 50 4590
rect 50 4538 230 4590
rect 230 4538 248 4590
rect 32 4536 248 4538
rect 1838 4898 1894 4906
rect 1838 4782 1840 4898
rect 1840 4782 1892 4898
rect 1892 4782 1894 4898
rect 1838 4772 1894 4782
rect 3306 7154 3362 7156
rect 3306 7100 3308 7154
rect 3308 7100 3362 7154
rect 3444 7100 3500 7156
rect 1170 4518 1226 4652
rect 2070 4338 2126 4474
rect 2758 4510 2814 4644
rect 2070 -23168 2126 -23158
rect 2070 -23284 2072 -23168
rect 2072 -23284 2124 -23168
rect 2124 -23284 2126 -23168
rect 2070 -23294 2126 -23284
<< metal3 >>
rect 2250 8016 2398 8020
rect -70 8014 3718 8016
rect -70 7958 2256 8014
rect 2392 7958 3718 8014
rect -70 7956 3718 7958
rect 2250 7952 2398 7956
rect 26 7860 254 7866
rect 26 7796 28 7860
rect 252 7796 254 7860
rect 26 7790 254 7796
rect 760 7676 908 7680
rect -70 7674 3718 7676
rect -70 7618 766 7674
rect 902 7618 3718 7674
rect -70 7616 3718 7618
rect 760 7612 908 7616
rect 8 7548 156 7554
rect 8 7476 14 7548
rect -70 7416 14 7476
rect 8 7412 14 7416
rect 150 7476 156 7548
rect 150 7416 3718 7476
rect 150 7412 156 7416
rect 8 7406 156 7412
rect 346 7316 574 7322
rect 346 7252 348 7316
rect 572 7252 574 7316
rect 346 7246 574 7252
rect 3300 7158 3368 7162
rect -70 7156 3368 7158
rect -70 7100 3306 7156
rect 3362 7100 3368 7156
rect -70 7098 3368 7100
rect 3300 7094 3368 7098
rect 3438 7160 3506 7162
rect 3438 7156 3718 7160
rect 3438 7100 3444 7156
rect 3500 7100 3718 7156
rect 3438 7094 3506 7100
rect 26 6772 254 6778
rect 26 6708 28 6772
rect 252 6708 254 6772
rect 26 6702 254 6708
rect 2 6536 70 6540
rect 1074 6536 1142 6540
rect 2 6534 1142 6536
rect 2 6478 8 6534
rect 64 6478 1080 6534
rect 1136 6478 1142 6534
rect 2 6476 1142 6478
rect 2 6472 70 6476
rect 1074 6472 1142 6476
rect 346 6228 574 6234
rect 346 6164 348 6228
rect 572 6164 574 6228
rect 346 6158 574 6164
rect 26 5684 254 5690
rect 26 5620 28 5684
rect 252 5620 254 5684
rect 26 5614 254 5620
rect 2 5446 70 5452
rect 2 5390 8 5446
rect 64 5444 70 5446
rect 1072 5444 1140 5448
rect 64 5442 1140 5444
rect 64 5390 1078 5442
rect 2 5386 1078 5390
rect 1134 5386 1140 5442
rect 2 5384 1140 5386
rect 1072 5380 1140 5384
rect 1544 5268 1550 5276
rect -8 5208 1550 5268
rect -8 4906 60 5208
rect 346 5140 574 5146
rect 346 5076 348 5140
rect 572 5076 574 5140
rect 1544 5132 1550 5208
rect 1614 5132 1620 5276
rect 346 5070 574 5076
rect -8 4772 -2 4906
rect 54 4772 60 4906
rect -8 4766 60 4772
rect 452 4906 520 4912
rect 1032 4906 1038 4912
rect 452 4772 458 4906
rect 514 4774 1038 4906
rect 514 4772 520 4774
rect 452 4766 520 4772
rect 1032 4768 1038 4774
rect 1102 4768 1108 4912
rect 1416 4768 1422 4912
rect 1486 4906 1900 4912
rect 1486 4772 1838 4906
rect 1894 4772 1900 4906
rect 1486 4768 1900 4772
rect 1832 4766 1900 4768
rect 1166 4658 1232 4662
rect 1164 4656 1232 4658
rect 26 4596 254 4602
rect 26 4532 28 4596
rect 252 4532 254 4596
rect 26 4526 254 4532
rect 1164 4512 1166 4656
rect 1230 4512 1232 4656
rect 1166 4506 1232 4512
rect 1294 4656 1360 4662
rect 1358 4608 1360 4656
rect 2752 4644 2820 4650
rect 2752 4608 2758 4644
rect 1358 4548 2758 4608
rect 1358 4512 1360 4548
rect 1294 4506 1360 4512
rect 2752 4510 2758 4548
rect 2814 4510 2820 4644
rect 2752 4504 2820 4510
rect 2064 4478 2132 4484
rect 2064 4334 2066 4478
rect 2130 4334 2132 4478
rect 2064 4328 2132 4334
rect 1032 -270 1038 -228
rect 952 -346 1038 -270
rect 1032 -372 1038 -346
rect 1102 -372 1108 -228
rect 1160 -4892 1166 -4850
rect 950 -4968 1166 -4892
rect 1160 -4994 1166 -4968
rect 1230 -4994 1236 -4850
rect 1288 -9514 1294 -9472
rect 950 -9590 1294 -9514
rect 1288 -9616 1294 -9590
rect 1358 -9616 1364 -9472
rect 1416 -14136 1422 -14094
rect 954 -14212 1422 -14136
rect 1416 -14238 1422 -14212
rect 1486 -14238 1492 -14094
rect 1544 -18758 1550 -18716
rect 952 -18834 1550 -18758
rect 1544 -18860 1550 -18834
rect 1614 -18860 1620 -18716
rect 2064 -23154 2132 -23152
rect 2060 -23298 2066 -23154
rect 2130 -23298 2136 -23154
rect 2064 -23300 2132 -23298
<< via3 >>
rect 28 7856 252 7860
rect 28 7800 32 7856
rect 32 7800 248 7856
rect 248 7800 252 7856
rect 28 7796 252 7800
rect 348 7312 572 7316
rect 348 7256 352 7312
rect 352 7256 568 7312
rect 568 7256 572 7312
rect 348 7252 572 7256
rect 28 6768 252 6772
rect 28 6712 32 6768
rect 32 6712 248 6768
rect 248 6712 252 6768
rect 28 6708 252 6712
rect 348 6224 572 6228
rect 348 6168 352 6224
rect 352 6168 568 6224
rect 568 6168 572 6224
rect 348 6164 572 6168
rect 28 5680 252 5684
rect 28 5624 70 5680
rect 70 5624 248 5680
rect 248 5624 252 5680
rect 28 5620 252 5624
rect 348 5136 572 5140
rect 348 5080 352 5136
rect 352 5080 568 5136
rect 568 5080 572 5136
rect 348 5076 572 5080
rect 1550 5132 1614 5276
rect 1038 4768 1102 4912
rect 1422 4768 1486 4912
rect 28 4592 252 4596
rect 28 4536 32 4592
rect 32 4536 248 4592
rect 248 4536 252 4592
rect 28 4532 252 4536
rect 1166 4652 1230 4656
rect 1166 4518 1170 4652
rect 1170 4518 1226 4652
rect 1226 4518 1230 4652
rect 1166 4512 1230 4518
rect 1294 4512 1358 4656
rect 2066 4474 2130 4478
rect 2066 4338 2070 4474
rect 2070 4338 2126 4474
rect 2126 4338 2130 4474
rect 2066 4334 2130 4338
rect 1038 -372 1102 -228
rect 1166 -4994 1230 -4850
rect 1294 -9616 1358 -9472
rect 1422 -14238 1486 -14094
rect 1550 -18860 1614 -18716
rect 2066 -23158 2130 -23154
rect 2066 -23294 2070 -23158
rect 2070 -23294 2126 -23158
rect 2126 -23294 2130 -23158
rect 2066 -23298 2130 -23294
<< metal4 >>
rect 26 7860 254 7862
rect 20 7796 28 7860
rect 252 7796 260 7860
rect 20 6772 260 7796
rect 20 6708 28 6772
rect 252 6708 260 6772
rect 20 5684 260 6708
rect 20 5620 28 5684
rect 252 5620 260 5684
rect 20 4596 260 5620
rect 20 4532 28 4596
rect 252 4532 260 4596
rect 20 -32354 260 4532
rect 340 7316 580 7860
rect 340 7252 348 7316
rect 572 7252 580 7316
rect 340 6228 580 7252
rect 340 6164 348 6228
rect 572 6164 580 6228
rect 340 5140 580 6164
rect 340 5076 348 5140
rect 572 5076 580 5140
rect 340 -32354 580 5076
rect 660 -32354 900 7860
rect 1548 5276 1616 5278
rect 1040 4914 1100 5156
rect 1036 4912 1104 4914
rect 1036 4768 1038 4912
rect 1102 4768 1104 4912
rect 1036 4766 1104 4768
rect 1040 -226 1100 4766
rect 1168 4658 1228 5156
rect 1296 4658 1356 5156
rect 1424 4914 1484 5156
rect 1548 5132 1550 5276
rect 1614 5132 1616 5276
rect 1548 5130 1616 5132
rect 1420 4912 1488 4914
rect 1420 4768 1422 4912
rect 1486 4768 1488 4912
rect 1420 4766 1488 4768
rect 1164 4656 1232 4658
rect 1164 4512 1166 4656
rect 1230 4512 1232 4656
rect 1164 4510 1232 4512
rect 1292 4656 1360 4658
rect 1292 4512 1294 4656
rect 1358 4512 1360 4656
rect 1292 4510 1360 4512
rect 1036 -228 1104 -226
rect 1036 -372 1038 -228
rect 1102 -372 1104 -228
rect 1036 -374 1104 -372
rect 1040 -23300 1100 -374
rect 1168 -4848 1228 4510
rect 1164 -4850 1232 -4848
rect 1164 -4994 1166 -4850
rect 1230 -4994 1232 -4850
rect 1164 -4996 1232 -4994
rect 1168 -23300 1228 -4996
rect 1296 -9470 1356 4510
rect 1292 -9472 1360 -9470
rect 1292 -9616 1294 -9472
rect 1358 -9616 1360 -9472
rect 1292 -9618 1360 -9616
rect 1296 -23300 1356 -9618
rect 1424 -14092 1484 4766
rect 1420 -14094 1488 -14092
rect 1420 -14238 1422 -14094
rect 1486 -14238 1488 -14094
rect 1420 -14240 1488 -14238
rect 1424 -23300 1484 -14240
rect 1552 -18714 1612 5130
rect 2068 4480 2128 4512
rect 2064 4478 2132 4480
rect 2064 4334 2066 4478
rect 2130 4334 2132 4478
rect 2064 4332 2132 4334
rect 1548 -18716 1616 -18714
rect 1548 -18860 1550 -18716
rect 1614 -18860 1616 -18716
rect 1548 -18862 1616 -18860
rect 1552 -23300 1612 -18862
rect 2068 -23152 2128 4332
rect 2064 -23154 2132 -23152
rect 2064 -23298 2066 -23154
rect 2130 -23298 2132 -23154
rect 2064 -23300 2132 -23298
use and  and_1
timestamp 1757283562
transform -1 0 444 0 -1 5110
box -38 -48 498 592
use and  and_2
timestamp 1757283562
transform -1 0 904 0 -1 5110
box -38 -48 498 592
use and  and_3
timestamp 1757283562
transform -1 0 1364 0 -1 5110
box -38 -48 498 592
use and  and_4
timestamp 1757283562
transform -1 0 1824 0 -1 5110
box -38 -48 498 592
use and  and_5
timestamp 1757283562
transform -1 0 2284 0 -1 5110
box -38 -48 498 592
use and  and_6
timestamp 1757283562
transform -1 0 2744 0 -1 5110
box -38 -48 498 592
use and  and_7
timestamp 1757283562
transform -1 0 3204 0 -1 5110
box -38 -48 498 592
use clkinv  clkinv_0
timestamp 1757283562
transform 1 0 76 0 1 7286
box -38 -48 314 592
use dff  dff_0
timestamp 1757283562
transform -1 0 1824 0 -1 7286
box -38 -48 1878 592
use dff  dff_1
timestamp 1757283562
transform 1 0 -16 0 1 6198
box -38 -48 1878 592
use dff  dff_3
timestamp 1757283562
transform -1 0 3664 0 -1 6198
box -38 -48 1878 592
use dff  dff_4
timestamp 1757283562
transform 1 0 1824 0 1 6198
box -38 -48 1878 592
use dff  dff_5
timestamp 1757283562
transform -1 0 3664 0 -1 7286
box -38 -48 1878 592
use dff  dff_6
timestamp 1757283562
transform -1 0 1824 0 -1 6198
box -38 -48 1878 592
use dff  dff_7
timestamp 1757283562
transform 1 0 -16 0 1 5110
box -38 -48 1878 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1675710598
transform -1 0 3296 0 -1 5110
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_1
timestamp 1675710598
transform -1 0 -16 0 -1 5110
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_2
timestamp 1675710598
transform -1 0 -16 0 -1 7286
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_3
timestamp 1675710598
transform -1 0 -16 0 -1 6198
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_4
timestamp 1675710598
transform 1 0 -108 0 1 7286
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_5
timestamp 1675710598
transform -1 0 3756 0 -1 7286
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_6
timestamp 1675710598
transform -1 0 3756 0 -1 6198
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_7
timestamp 1675710598
transform 1 0 -108 0 1 5110
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_8
timestamp 1675710598
transform 1 0 -108 0 1 6198
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_9
timestamp 1675710598
transform 1 0 3664 0 1 6198
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_10
timestamp 1675710598
transform 1 0 3664 0 1 5110
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_11
timestamp 1675710598
transform -1 0 3756 0 -1 5110
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_12
timestamp 1675710598
transform -1 0 3664 0 -1 5110
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_13
timestamp 1675710598
transform -1 0 3572 0 -1 5110
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_14
timestamp 1675710598
transform -1 0 3480 0 -1 5110
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_15
timestamp 1675710598
transform -1 0 3388 0 -1 5110
box -38 -48 130 592
use tt_asw_3v3  tt_asw_3v3_0
timestamp 1757283562
transform 1 0 0 0 1 -23110
box 0 0 3612 4352
use tt_asw_3v3  tt_asw_3v3_1
timestamp 1757283562
transform 1 0 0 0 1 0
box 0 0 3612 4352
use tt_asw_3v3  tt_asw_3v3_2
timestamp 1757283562
transform 1 0 0 0 1 -4622
box 0 0 3612 4352
use tt_asw_3v3  tt_asw_3v3_3
timestamp 1757283562
transform 1 0 0 0 1 -9244
box 0 0 3612 4352
use tt_asw_3v3  tt_asw_3v3_4
timestamp 1757283562
transform 1 0 0 0 1 -13866
box 0 0 3612 4352
use tt_asw_3v3  tt_asw_3v3_5
timestamp 1757283562
transform 1 0 0 0 1 -18488
box 0 0 3612 4352
use tt_asw_3v3  tt_asw_3v3_7
timestamp 1757283562
transform 1 0 0 0 1 -27732
box 0 0 3612 4352
<< labels >>
flabel locali s 1853 4855 1887 4889 0 FreeSans 250 180 0 0 X
port 7 nsew signal output
flabel locali s 1853 4787 1887 4821 0 FreeSans 250 180 0 0 X
port 7 nsew signal output
<< end >>
