magic
tech sky130A
magscale 1 2
timestamp 1757105855
<< error_p >>
rect -101 -174 -100 174
rect 100 -174 101 174
<< nwell >>
rect -3196 -3269 3196 3269
<< mvpmos >>
rect -2938 1972 -2738 2972
rect -2680 1972 -2480 2972
rect -2422 1972 -2222 2972
rect -2164 1972 -1964 2972
rect -1906 1972 -1706 2972
rect -1648 1972 -1448 2972
rect -1390 1972 -1190 2972
rect -1132 1972 -932 2972
rect -874 1972 -674 2972
rect -616 1972 -416 2972
rect -358 1972 -158 2972
rect -100 1972 100 2972
rect 158 1972 358 2972
rect 416 1972 616 2972
rect 674 1972 874 2972
rect 932 1972 1132 2972
rect 1190 1972 1390 2972
rect 1448 1972 1648 2972
rect 1706 1972 1906 2972
rect 1964 1972 2164 2972
rect 2222 1972 2422 2972
rect 2480 1972 2680 2972
rect 2738 1972 2938 2972
rect -2938 736 -2738 1736
rect -2680 736 -2480 1736
rect -2422 736 -2222 1736
rect -2164 736 -1964 1736
rect -1906 736 -1706 1736
rect -1648 736 -1448 1736
rect -1390 736 -1190 1736
rect -1132 736 -932 1736
rect -874 736 -674 1736
rect -616 736 -416 1736
rect -358 736 -158 1736
rect -100 736 100 1736
rect 158 736 358 1736
rect 416 736 616 1736
rect 674 736 874 1736
rect 932 736 1132 1736
rect 1190 736 1390 1736
rect 1448 736 1648 1736
rect 1706 736 1906 1736
rect 1964 736 2164 1736
rect 2222 736 2422 1736
rect 2480 736 2680 1736
rect 2738 736 2938 1736
rect -2938 -500 -2738 500
rect -2680 -500 -2480 500
rect -2422 -500 -2222 500
rect -2164 -500 -1964 500
rect -1906 -500 -1706 500
rect -1648 -500 -1448 500
rect -1390 -500 -1190 500
rect -1132 -500 -932 500
rect -874 -500 -674 500
rect -616 -500 -416 500
rect -358 -500 -158 500
rect -100 -500 100 500
rect 158 -500 358 500
rect 416 -500 616 500
rect 674 -500 874 500
rect 932 -500 1132 500
rect 1190 -500 1390 500
rect 1448 -500 1648 500
rect 1706 -500 1906 500
rect 1964 -500 2164 500
rect 2222 -500 2422 500
rect 2480 -500 2680 500
rect 2738 -500 2938 500
rect -2938 -1736 -2738 -736
rect -2680 -1736 -2480 -736
rect -2422 -1736 -2222 -736
rect -2164 -1736 -1964 -736
rect -1906 -1736 -1706 -736
rect -1648 -1736 -1448 -736
rect -1390 -1736 -1190 -736
rect -1132 -1736 -932 -736
rect -874 -1736 -674 -736
rect -616 -1736 -416 -736
rect -358 -1736 -158 -736
rect -100 -1736 100 -736
rect 158 -1736 358 -736
rect 416 -1736 616 -736
rect 674 -1736 874 -736
rect 932 -1736 1132 -736
rect 1190 -1736 1390 -736
rect 1448 -1736 1648 -736
rect 1706 -1736 1906 -736
rect 1964 -1736 2164 -736
rect 2222 -1736 2422 -736
rect 2480 -1736 2680 -736
rect 2738 -1736 2938 -736
rect -2938 -2972 -2738 -1972
rect -2680 -2972 -2480 -1972
rect -2422 -2972 -2222 -1972
rect -2164 -2972 -1964 -1972
rect -1906 -2972 -1706 -1972
rect -1648 -2972 -1448 -1972
rect -1390 -2972 -1190 -1972
rect -1132 -2972 -932 -1972
rect -874 -2972 -674 -1972
rect -616 -2972 -416 -1972
rect -358 -2972 -158 -1972
rect -100 -2972 100 -1972
rect 158 -2972 358 -1972
rect 416 -2972 616 -1972
rect 674 -2972 874 -1972
rect 932 -2972 1132 -1972
rect 1190 -2972 1390 -1972
rect 1448 -2972 1648 -1972
rect 1706 -2972 1906 -1972
rect 1964 -2972 2164 -1972
rect 2222 -2972 2422 -1972
rect 2480 -2972 2680 -1972
rect 2738 -2972 2938 -1972
<< mvpdiff >>
rect -2996 2960 -2938 2972
rect -2996 1984 -2984 2960
rect -2950 1984 -2938 2960
rect -2996 1972 -2938 1984
rect -2738 2960 -2680 2972
rect -2738 1984 -2726 2960
rect -2692 1984 -2680 2960
rect -2738 1972 -2680 1984
rect -2480 2960 -2422 2972
rect -2480 1984 -2468 2960
rect -2434 1984 -2422 2960
rect -2480 1972 -2422 1984
rect -2222 2960 -2164 2972
rect -2222 1984 -2210 2960
rect -2176 1984 -2164 2960
rect -2222 1972 -2164 1984
rect -1964 2960 -1906 2972
rect -1964 1984 -1952 2960
rect -1918 1984 -1906 2960
rect -1964 1972 -1906 1984
rect -1706 2960 -1648 2972
rect -1706 1984 -1694 2960
rect -1660 1984 -1648 2960
rect -1706 1972 -1648 1984
rect -1448 2960 -1390 2972
rect -1448 1984 -1436 2960
rect -1402 1984 -1390 2960
rect -1448 1972 -1390 1984
rect -1190 2960 -1132 2972
rect -1190 1984 -1178 2960
rect -1144 1984 -1132 2960
rect -1190 1972 -1132 1984
rect -932 2960 -874 2972
rect -932 1984 -920 2960
rect -886 1984 -874 2960
rect -932 1972 -874 1984
rect -674 2960 -616 2972
rect -674 1984 -662 2960
rect -628 1984 -616 2960
rect -674 1972 -616 1984
rect -416 2960 -358 2972
rect -416 1984 -404 2960
rect -370 1984 -358 2960
rect -416 1972 -358 1984
rect -158 2960 -100 2972
rect -158 1984 -146 2960
rect -112 1984 -100 2960
rect -158 1972 -100 1984
rect 100 2960 158 2972
rect 100 1984 112 2960
rect 146 1984 158 2960
rect 100 1972 158 1984
rect 358 2960 416 2972
rect 358 1984 370 2960
rect 404 1984 416 2960
rect 358 1972 416 1984
rect 616 2960 674 2972
rect 616 1984 628 2960
rect 662 1984 674 2960
rect 616 1972 674 1984
rect 874 2960 932 2972
rect 874 1984 886 2960
rect 920 1984 932 2960
rect 874 1972 932 1984
rect 1132 2960 1190 2972
rect 1132 1984 1144 2960
rect 1178 1984 1190 2960
rect 1132 1972 1190 1984
rect 1390 2960 1448 2972
rect 1390 1984 1402 2960
rect 1436 1984 1448 2960
rect 1390 1972 1448 1984
rect 1648 2960 1706 2972
rect 1648 1984 1660 2960
rect 1694 1984 1706 2960
rect 1648 1972 1706 1984
rect 1906 2960 1964 2972
rect 1906 1984 1918 2960
rect 1952 1984 1964 2960
rect 1906 1972 1964 1984
rect 2164 2960 2222 2972
rect 2164 1984 2176 2960
rect 2210 1984 2222 2960
rect 2164 1972 2222 1984
rect 2422 2960 2480 2972
rect 2422 1984 2434 2960
rect 2468 1984 2480 2960
rect 2422 1972 2480 1984
rect 2680 2960 2738 2972
rect 2680 1984 2692 2960
rect 2726 1984 2738 2960
rect 2680 1972 2738 1984
rect 2938 2960 2996 2972
rect 2938 1984 2950 2960
rect 2984 1984 2996 2960
rect 2938 1972 2996 1984
rect -2996 1724 -2938 1736
rect -2996 748 -2984 1724
rect -2950 748 -2938 1724
rect -2996 736 -2938 748
rect -2738 1724 -2680 1736
rect -2738 748 -2726 1724
rect -2692 748 -2680 1724
rect -2738 736 -2680 748
rect -2480 1724 -2422 1736
rect -2480 748 -2468 1724
rect -2434 748 -2422 1724
rect -2480 736 -2422 748
rect -2222 1724 -2164 1736
rect -2222 748 -2210 1724
rect -2176 748 -2164 1724
rect -2222 736 -2164 748
rect -1964 1724 -1906 1736
rect -1964 748 -1952 1724
rect -1918 748 -1906 1724
rect -1964 736 -1906 748
rect -1706 1724 -1648 1736
rect -1706 748 -1694 1724
rect -1660 748 -1648 1724
rect -1706 736 -1648 748
rect -1448 1724 -1390 1736
rect -1448 748 -1436 1724
rect -1402 748 -1390 1724
rect -1448 736 -1390 748
rect -1190 1724 -1132 1736
rect -1190 748 -1178 1724
rect -1144 748 -1132 1724
rect -1190 736 -1132 748
rect -932 1724 -874 1736
rect -932 748 -920 1724
rect -886 748 -874 1724
rect -932 736 -874 748
rect -674 1724 -616 1736
rect -674 748 -662 1724
rect -628 748 -616 1724
rect -674 736 -616 748
rect -416 1724 -358 1736
rect -416 748 -404 1724
rect -370 748 -358 1724
rect -416 736 -358 748
rect -158 1724 -100 1736
rect -158 748 -146 1724
rect -112 748 -100 1724
rect -158 736 -100 748
rect 100 1724 158 1736
rect 100 748 112 1724
rect 146 748 158 1724
rect 100 736 158 748
rect 358 1724 416 1736
rect 358 748 370 1724
rect 404 748 416 1724
rect 358 736 416 748
rect 616 1724 674 1736
rect 616 748 628 1724
rect 662 748 674 1724
rect 616 736 674 748
rect 874 1724 932 1736
rect 874 748 886 1724
rect 920 748 932 1724
rect 874 736 932 748
rect 1132 1724 1190 1736
rect 1132 748 1144 1724
rect 1178 748 1190 1724
rect 1132 736 1190 748
rect 1390 1724 1448 1736
rect 1390 748 1402 1724
rect 1436 748 1448 1724
rect 1390 736 1448 748
rect 1648 1724 1706 1736
rect 1648 748 1660 1724
rect 1694 748 1706 1724
rect 1648 736 1706 748
rect 1906 1724 1964 1736
rect 1906 748 1918 1724
rect 1952 748 1964 1724
rect 1906 736 1964 748
rect 2164 1724 2222 1736
rect 2164 748 2176 1724
rect 2210 748 2222 1724
rect 2164 736 2222 748
rect 2422 1724 2480 1736
rect 2422 748 2434 1724
rect 2468 748 2480 1724
rect 2422 736 2480 748
rect 2680 1724 2738 1736
rect 2680 748 2692 1724
rect 2726 748 2738 1724
rect 2680 736 2738 748
rect 2938 1724 2996 1736
rect 2938 748 2950 1724
rect 2984 748 2996 1724
rect 2938 736 2996 748
rect -2996 488 -2938 500
rect -2996 -488 -2984 488
rect -2950 -488 -2938 488
rect -2996 -500 -2938 -488
rect -2738 488 -2680 500
rect -2738 -488 -2726 488
rect -2692 -488 -2680 488
rect -2738 -500 -2680 -488
rect -2480 488 -2422 500
rect -2480 -488 -2468 488
rect -2434 -488 -2422 488
rect -2480 -500 -2422 -488
rect -2222 488 -2164 500
rect -2222 -488 -2210 488
rect -2176 -488 -2164 488
rect -2222 -500 -2164 -488
rect -1964 488 -1906 500
rect -1964 -488 -1952 488
rect -1918 -488 -1906 488
rect -1964 -500 -1906 -488
rect -1706 488 -1648 500
rect -1706 -488 -1694 488
rect -1660 -488 -1648 488
rect -1706 -500 -1648 -488
rect -1448 488 -1390 500
rect -1448 -488 -1436 488
rect -1402 -488 -1390 488
rect -1448 -500 -1390 -488
rect -1190 488 -1132 500
rect -1190 -488 -1178 488
rect -1144 -488 -1132 488
rect -1190 -500 -1132 -488
rect -932 488 -874 500
rect -932 -488 -920 488
rect -886 -488 -874 488
rect -932 -500 -874 -488
rect -674 488 -616 500
rect -674 -488 -662 488
rect -628 -488 -616 488
rect -674 -500 -616 -488
rect -416 488 -358 500
rect -416 -488 -404 488
rect -370 -488 -358 488
rect -416 -500 -358 -488
rect -158 488 -100 500
rect -158 -488 -146 488
rect -112 -488 -100 488
rect -158 -500 -100 -488
rect 100 488 158 500
rect 100 -488 112 488
rect 146 -488 158 488
rect 100 -500 158 -488
rect 358 488 416 500
rect 358 -488 370 488
rect 404 -488 416 488
rect 358 -500 416 -488
rect 616 488 674 500
rect 616 -488 628 488
rect 662 -488 674 488
rect 616 -500 674 -488
rect 874 488 932 500
rect 874 -488 886 488
rect 920 -488 932 488
rect 874 -500 932 -488
rect 1132 488 1190 500
rect 1132 -488 1144 488
rect 1178 -488 1190 488
rect 1132 -500 1190 -488
rect 1390 488 1448 500
rect 1390 -488 1402 488
rect 1436 -488 1448 488
rect 1390 -500 1448 -488
rect 1648 488 1706 500
rect 1648 -488 1660 488
rect 1694 -488 1706 488
rect 1648 -500 1706 -488
rect 1906 488 1964 500
rect 1906 -488 1918 488
rect 1952 -488 1964 488
rect 1906 -500 1964 -488
rect 2164 488 2222 500
rect 2164 -488 2176 488
rect 2210 -488 2222 488
rect 2164 -500 2222 -488
rect 2422 488 2480 500
rect 2422 -488 2434 488
rect 2468 -488 2480 488
rect 2422 -500 2480 -488
rect 2680 488 2738 500
rect 2680 -488 2692 488
rect 2726 -488 2738 488
rect 2680 -500 2738 -488
rect 2938 488 2996 500
rect 2938 -488 2950 488
rect 2984 -488 2996 488
rect 2938 -500 2996 -488
rect -2996 -748 -2938 -736
rect -2996 -1724 -2984 -748
rect -2950 -1724 -2938 -748
rect -2996 -1736 -2938 -1724
rect -2738 -748 -2680 -736
rect -2738 -1724 -2726 -748
rect -2692 -1724 -2680 -748
rect -2738 -1736 -2680 -1724
rect -2480 -748 -2422 -736
rect -2480 -1724 -2468 -748
rect -2434 -1724 -2422 -748
rect -2480 -1736 -2422 -1724
rect -2222 -748 -2164 -736
rect -2222 -1724 -2210 -748
rect -2176 -1724 -2164 -748
rect -2222 -1736 -2164 -1724
rect -1964 -748 -1906 -736
rect -1964 -1724 -1952 -748
rect -1918 -1724 -1906 -748
rect -1964 -1736 -1906 -1724
rect -1706 -748 -1648 -736
rect -1706 -1724 -1694 -748
rect -1660 -1724 -1648 -748
rect -1706 -1736 -1648 -1724
rect -1448 -748 -1390 -736
rect -1448 -1724 -1436 -748
rect -1402 -1724 -1390 -748
rect -1448 -1736 -1390 -1724
rect -1190 -748 -1132 -736
rect -1190 -1724 -1178 -748
rect -1144 -1724 -1132 -748
rect -1190 -1736 -1132 -1724
rect -932 -748 -874 -736
rect -932 -1724 -920 -748
rect -886 -1724 -874 -748
rect -932 -1736 -874 -1724
rect -674 -748 -616 -736
rect -674 -1724 -662 -748
rect -628 -1724 -616 -748
rect -674 -1736 -616 -1724
rect -416 -748 -358 -736
rect -416 -1724 -404 -748
rect -370 -1724 -358 -748
rect -416 -1736 -358 -1724
rect -158 -748 -100 -736
rect -158 -1724 -146 -748
rect -112 -1724 -100 -748
rect -158 -1736 -100 -1724
rect 100 -748 158 -736
rect 100 -1724 112 -748
rect 146 -1724 158 -748
rect 100 -1736 158 -1724
rect 358 -748 416 -736
rect 358 -1724 370 -748
rect 404 -1724 416 -748
rect 358 -1736 416 -1724
rect 616 -748 674 -736
rect 616 -1724 628 -748
rect 662 -1724 674 -748
rect 616 -1736 674 -1724
rect 874 -748 932 -736
rect 874 -1724 886 -748
rect 920 -1724 932 -748
rect 874 -1736 932 -1724
rect 1132 -748 1190 -736
rect 1132 -1724 1144 -748
rect 1178 -1724 1190 -748
rect 1132 -1736 1190 -1724
rect 1390 -748 1448 -736
rect 1390 -1724 1402 -748
rect 1436 -1724 1448 -748
rect 1390 -1736 1448 -1724
rect 1648 -748 1706 -736
rect 1648 -1724 1660 -748
rect 1694 -1724 1706 -748
rect 1648 -1736 1706 -1724
rect 1906 -748 1964 -736
rect 1906 -1724 1918 -748
rect 1952 -1724 1964 -748
rect 1906 -1736 1964 -1724
rect 2164 -748 2222 -736
rect 2164 -1724 2176 -748
rect 2210 -1724 2222 -748
rect 2164 -1736 2222 -1724
rect 2422 -748 2480 -736
rect 2422 -1724 2434 -748
rect 2468 -1724 2480 -748
rect 2422 -1736 2480 -1724
rect 2680 -748 2738 -736
rect 2680 -1724 2692 -748
rect 2726 -1724 2738 -748
rect 2680 -1736 2738 -1724
rect 2938 -748 2996 -736
rect 2938 -1724 2950 -748
rect 2984 -1724 2996 -748
rect 2938 -1736 2996 -1724
rect -2996 -1984 -2938 -1972
rect -2996 -2960 -2984 -1984
rect -2950 -2960 -2938 -1984
rect -2996 -2972 -2938 -2960
rect -2738 -1984 -2680 -1972
rect -2738 -2960 -2726 -1984
rect -2692 -2960 -2680 -1984
rect -2738 -2972 -2680 -2960
rect -2480 -1984 -2422 -1972
rect -2480 -2960 -2468 -1984
rect -2434 -2960 -2422 -1984
rect -2480 -2972 -2422 -2960
rect -2222 -1984 -2164 -1972
rect -2222 -2960 -2210 -1984
rect -2176 -2960 -2164 -1984
rect -2222 -2972 -2164 -2960
rect -1964 -1984 -1906 -1972
rect -1964 -2960 -1952 -1984
rect -1918 -2960 -1906 -1984
rect -1964 -2972 -1906 -2960
rect -1706 -1984 -1648 -1972
rect -1706 -2960 -1694 -1984
rect -1660 -2960 -1648 -1984
rect -1706 -2972 -1648 -2960
rect -1448 -1984 -1390 -1972
rect -1448 -2960 -1436 -1984
rect -1402 -2960 -1390 -1984
rect -1448 -2972 -1390 -2960
rect -1190 -1984 -1132 -1972
rect -1190 -2960 -1178 -1984
rect -1144 -2960 -1132 -1984
rect -1190 -2972 -1132 -2960
rect -932 -1984 -874 -1972
rect -932 -2960 -920 -1984
rect -886 -2960 -874 -1984
rect -932 -2972 -874 -2960
rect -674 -1984 -616 -1972
rect -674 -2960 -662 -1984
rect -628 -2960 -616 -1984
rect -674 -2972 -616 -2960
rect -416 -1984 -358 -1972
rect -416 -2960 -404 -1984
rect -370 -2960 -358 -1984
rect -416 -2972 -358 -2960
rect -158 -1984 -100 -1972
rect -158 -2960 -146 -1984
rect -112 -2960 -100 -1984
rect -158 -2972 -100 -2960
rect 100 -1984 158 -1972
rect 100 -2960 112 -1984
rect 146 -2960 158 -1984
rect 100 -2972 158 -2960
rect 358 -1984 416 -1972
rect 358 -2960 370 -1984
rect 404 -2960 416 -1984
rect 358 -2972 416 -2960
rect 616 -1984 674 -1972
rect 616 -2960 628 -1984
rect 662 -2960 674 -1984
rect 616 -2972 674 -2960
rect 874 -1984 932 -1972
rect 874 -2960 886 -1984
rect 920 -2960 932 -1984
rect 874 -2972 932 -2960
rect 1132 -1984 1190 -1972
rect 1132 -2960 1144 -1984
rect 1178 -2960 1190 -1984
rect 1132 -2972 1190 -2960
rect 1390 -1984 1448 -1972
rect 1390 -2960 1402 -1984
rect 1436 -2960 1448 -1984
rect 1390 -2972 1448 -2960
rect 1648 -1984 1706 -1972
rect 1648 -2960 1660 -1984
rect 1694 -2960 1706 -1984
rect 1648 -2972 1706 -2960
rect 1906 -1984 1964 -1972
rect 1906 -2960 1918 -1984
rect 1952 -2960 1964 -1984
rect 1906 -2972 1964 -2960
rect 2164 -1984 2222 -1972
rect 2164 -2960 2176 -1984
rect 2210 -2960 2222 -1984
rect 2164 -2972 2222 -2960
rect 2422 -1984 2480 -1972
rect 2422 -2960 2434 -1984
rect 2468 -2960 2480 -1984
rect 2422 -2972 2480 -2960
rect 2680 -1984 2738 -1972
rect 2680 -2960 2692 -1984
rect 2726 -2960 2738 -1984
rect 2680 -2972 2738 -2960
rect 2938 -1984 2996 -1972
rect 2938 -2960 2950 -1984
rect 2984 -2960 2996 -1984
rect 2938 -2972 2996 -2960
<< mvpdiffc >>
rect -2984 1984 -2950 2960
rect -2726 1984 -2692 2960
rect -2468 1984 -2434 2960
rect -2210 1984 -2176 2960
rect -1952 1984 -1918 2960
rect -1694 1984 -1660 2960
rect -1436 1984 -1402 2960
rect -1178 1984 -1144 2960
rect -920 1984 -886 2960
rect -662 1984 -628 2960
rect -404 1984 -370 2960
rect -146 1984 -112 2960
rect 112 1984 146 2960
rect 370 1984 404 2960
rect 628 1984 662 2960
rect 886 1984 920 2960
rect 1144 1984 1178 2960
rect 1402 1984 1436 2960
rect 1660 1984 1694 2960
rect 1918 1984 1952 2960
rect 2176 1984 2210 2960
rect 2434 1984 2468 2960
rect 2692 1984 2726 2960
rect 2950 1984 2984 2960
rect -2984 748 -2950 1724
rect -2726 748 -2692 1724
rect -2468 748 -2434 1724
rect -2210 748 -2176 1724
rect -1952 748 -1918 1724
rect -1694 748 -1660 1724
rect -1436 748 -1402 1724
rect -1178 748 -1144 1724
rect -920 748 -886 1724
rect -662 748 -628 1724
rect -404 748 -370 1724
rect -146 748 -112 1724
rect 112 748 146 1724
rect 370 748 404 1724
rect 628 748 662 1724
rect 886 748 920 1724
rect 1144 748 1178 1724
rect 1402 748 1436 1724
rect 1660 748 1694 1724
rect 1918 748 1952 1724
rect 2176 748 2210 1724
rect 2434 748 2468 1724
rect 2692 748 2726 1724
rect 2950 748 2984 1724
rect -2984 -488 -2950 488
rect -2726 -488 -2692 488
rect -2468 -488 -2434 488
rect -2210 -488 -2176 488
rect -1952 -488 -1918 488
rect -1694 -488 -1660 488
rect -1436 -488 -1402 488
rect -1178 -488 -1144 488
rect -920 -488 -886 488
rect -662 -488 -628 488
rect -404 -488 -370 488
rect -146 -488 -112 488
rect 112 -488 146 488
rect 370 -488 404 488
rect 628 -488 662 488
rect 886 -488 920 488
rect 1144 -488 1178 488
rect 1402 -488 1436 488
rect 1660 -488 1694 488
rect 1918 -488 1952 488
rect 2176 -488 2210 488
rect 2434 -488 2468 488
rect 2692 -488 2726 488
rect 2950 -488 2984 488
rect -2984 -1724 -2950 -748
rect -2726 -1724 -2692 -748
rect -2468 -1724 -2434 -748
rect -2210 -1724 -2176 -748
rect -1952 -1724 -1918 -748
rect -1694 -1724 -1660 -748
rect -1436 -1724 -1402 -748
rect -1178 -1724 -1144 -748
rect -920 -1724 -886 -748
rect -662 -1724 -628 -748
rect -404 -1724 -370 -748
rect -146 -1724 -112 -748
rect 112 -1724 146 -748
rect 370 -1724 404 -748
rect 628 -1724 662 -748
rect 886 -1724 920 -748
rect 1144 -1724 1178 -748
rect 1402 -1724 1436 -748
rect 1660 -1724 1694 -748
rect 1918 -1724 1952 -748
rect 2176 -1724 2210 -748
rect 2434 -1724 2468 -748
rect 2692 -1724 2726 -748
rect 2950 -1724 2984 -748
rect -2984 -2960 -2950 -1984
rect -2726 -2960 -2692 -1984
rect -2468 -2960 -2434 -1984
rect -2210 -2960 -2176 -1984
rect -1952 -2960 -1918 -1984
rect -1694 -2960 -1660 -1984
rect -1436 -2960 -1402 -1984
rect -1178 -2960 -1144 -1984
rect -920 -2960 -886 -1984
rect -662 -2960 -628 -1984
rect -404 -2960 -370 -1984
rect -146 -2960 -112 -1984
rect 112 -2960 146 -1984
rect 370 -2960 404 -1984
rect 628 -2960 662 -1984
rect 886 -2960 920 -1984
rect 1144 -2960 1178 -1984
rect 1402 -2960 1436 -1984
rect 1660 -2960 1694 -1984
rect 1918 -2960 1952 -1984
rect 2176 -2960 2210 -1984
rect 2434 -2960 2468 -1984
rect 2692 -2960 2726 -1984
rect 2950 -2960 2984 -1984
<< mvnsubdiff >>
rect -3130 3191 3130 3203
rect -3130 3157 -3022 3191
rect 3022 3157 3130 3191
rect -3130 3145 3130 3157
rect -3130 3095 -3072 3145
rect -3130 -3095 -3118 3095
rect -3084 -3095 -3072 3095
rect 3072 3095 3130 3145
rect -3130 -3145 -3072 -3095
rect 3072 -3095 3084 3095
rect 3118 -3095 3130 3095
rect 3072 -3145 3130 -3095
rect -3130 -3157 3130 -3145
rect -3130 -3191 -3022 -3157
rect 3022 -3191 3130 -3157
rect -3130 -3203 3130 -3191
<< mvnsubdiffcont >>
rect -3022 3157 3022 3191
rect -3118 -3095 -3084 3095
rect 3084 -3095 3118 3095
rect -3022 -3191 3022 -3157
<< poly >>
rect -2938 3053 -2738 3069
rect -2938 3019 -2922 3053
rect -2754 3019 -2738 3053
rect -2938 2972 -2738 3019
rect -2680 3053 -2480 3069
rect -2680 3019 -2664 3053
rect -2496 3019 -2480 3053
rect -2680 2972 -2480 3019
rect -2422 3053 -2222 3069
rect -2422 3019 -2406 3053
rect -2238 3019 -2222 3053
rect -2422 2972 -2222 3019
rect -2164 3053 -1964 3069
rect -2164 3019 -2148 3053
rect -1980 3019 -1964 3053
rect -2164 2972 -1964 3019
rect -1906 3053 -1706 3069
rect -1906 3019 -1890 3053
rect -1722 3019 -1706 3053
rect -1906 2972 -1706 3019
rect -1648 3053 -1448 3069
rect -1648 3019 -1632 3053
rect -1464 3019 -1448 3053
rect -1648 2972 -1448 3019
rect -1390 3053 -1190 3069
rect -1390 3019 -1374 3053
rect -1206 3019 -1190 3053
rect -1390 2972 -1190 3019
rect -1132 3053 -932 3069
rect -1132 3019 -1116 3053
rect -948 3019 -932 3053
rect -1132 2972 -932 3019
rect -874 3053 -674 3069
rect -874 3019 -858 3053
rect -690 3019 -674 3053
rect -874 2972 -674 3019
rect -616 3053 -416 3069
rect -616 3019 -600 3053
rect -432 3019 -416 3053
rect -616 2972 -416 3019
rect -358 3053 -158 3069
rect -358 3019 -342 3053
rect -174 3019 -158 3053
rect -358 2972 -158 3019
rect -100 3053 100 3069
rect -100 3019 -84 3053
rect 84 3019 100 3053
rect -100 2972 100 3019
rect 158 3053 358 3069
rect 158 3019 174 3053
rect 342 3019 358 3053
rect 158 2972 358 3019
rect 416 3053 616 3069
rect 416 3019 432 3053
rect 600 3019 616 3053
rect 416 2972 616 3019
rect 674 3053 874 3069
rect 674 3019 690 3053
rect 858 3019 874 3053
rect 674 2972 874 3019
rect 932 3053 1132 3069
rect 932 3019 948 3053
rect 1116 3019 1132 3053
rect 932 2972 1132 3019
rect 1190 3053 1390 3069
rect 1190 3019 1206 3053
rect 1374 3019 1390 3053
rect 1190 2972 1390 3019
rect 1448 3053 1648 3069
rect 1448 3019 1464 3053
rect 1632 3019 1648 3053
rect 1448 2972 1648 3019
rect 1706 3053 1906 3069
rect 1706 3019 1722 3053
rect 1890 3019 1906 3053
rect 1706 2972 1906 3019
rect 1964 3053 2164 3069
rect 1964 3019 1980 3053
rect 2148 3019 2164 3053
rect 1964 2972 2164 3019
rect 2222 3053 2422 3069
rect 2222 3019 2238 3053
rect 2406 3019 2422 3053
rect 2222 2972 2422 3019
rect 2480 3053 2680 3069
rect 2480 3019 2496 3053
rect 2664 3019 2680 3053
rect 2480 2972 2680 3019
rect 2738 3053 2938 3069
rect 2738 3019 2754 3053
rect 2922 3019 2938 3053
rect 2738 2972 2938 3019
rect -2938 1925 -2738 1972
rect -2938 1891 -2922 1925
rect -2754 1891 -2738 1925
rect -2938 1875 -2738 1891
rect -2680 1925 -2480 1972
rect -2680 1891 -2664 1925
rect -2496 1891 -2480 1925
rect -2680 1875 -2480 1891
rect -2422 1925 -2222 1972
rect -2422 1891 -2406 1925
rect -2238 1891 -2222 1925
rect -2422 1875 -2222 1891
rect -2164 1925 -1964 1972
rect -2164 1891 -2148 1925
rect -1980 1891 -1964 1925
rect -2164 1875 -1964 1891
rect -1906 1925 -1706 1972
rect -1906 1891 -1890 1925
rect -1722 1891 -1706 1925
rect -1906 1875 -1706 1891
rect -1648 1925 -1448 1972
rect -1648 1891 -1632 1925
rect -1464 1891 -1448 1925
rect -1648 1875 -1448 1891
rect -1390 1925 -1190 1972
rect -1390 1891 -1374 1925
rect -1206 1891 -1190 1925
rect -1390 1875 -1190 1891
rect -1132 1925 -932 1972
rect -1132 1891 -1116 1925
rect -948 1891 -932 1925
rect -1132 1875 -932 1891
rect -874 1925 -674 1972
rect -874 1891 -858 1925
rect -690 1891 -674 1925
rect -874 1875 -674 1891
rect -616 1925 -416 1972
rect -616 1891 -600 1925
rect -432 1891 -416 1925
rect -616 1875 -416 1891
rect -358 1925 -158 1972
rect -358 1891 -342 1925
rect -174 1891 -158 1925
rect -358 1875 -158 1891
rect -100 1925 100 1972
rect -100 1891 -84 1925
rect 84 1891 100 1925
rect -100 1875 100 1891
rect 158 1925 358 1972
rect 158 1891 174 1925
rect 342 1891 358 1925
rect 158 1875 358 1891
rect 416 1925 616 1972
rect 416 1891 432 1925
rect 600 1891 616 1925
rect 416 1875 616 1891
rect 674 1925 874 1972
rect 674 1891 690 1925
rect 858 1891 874 1925
rect 674 1875 874 1891
rect 932 1925 1132 1972
rect 932 1891 948 1925
rect 1116 1891 1132 1925
rect 932 1875 1132 1891
rect 1190 1925 1390 1972
rect 1190 1891 1206 1925
rect 1374 1891 1390 1925
rect 1190 1875 1390 1891
rect 1448 1925 1648 1972
rect 1448 1891 1464 1925
rect 1632 1891 1648 1925
rect 1448 1875 1648 1891
rect 1706 1925 1906 1972
rect 1706 1891 1722 1925
rect 1890 1891 1906 1925
rect 1706 1875 1906 1891
rect 1964 1925 2164 1972
rect 1964 1891 1980 1925
rect 2148 1891 2164 1925
rect 1964 1875 2164 1891
rect 2222 1925 2422 1972
rect 2222 1891 2238 1925
rect 2406 1891 2422 1925
rect 2222 1875 2422 1891
rect 2480 1925 2680 1972
rect 2480 1891 2496 1925
rect 2664 1891 2680 1925
rect 2480 1875 2680 1891
rect 2738 1925 2938 1972
rect 2738 1891 2754 1925
rect 2922 1891 2938 1925
rect 2738 1875 2938 1891
rect -2938 1817 -2738 1833
rect -2938 1783 -2922 1817
rect -2754 1783 -2738 1817
rect -2938 1736 -2738 1783
rect -2680 1817 -2480 1833
rect -2680 1783 -2664 1817
rect -2496 1783 -2480 1817
rect -2680 1736 -2480 1783
rect -2422 1817 -2222 1833
rect -2422 1783 -2406 1817
rect -2238 1783 -2222 1817
rect -2422 1736 -2222 1783
rect -2164 1817 -1964 1833
rect -2164 1783 -2148 1817
rect -1980 1783 -1964 1817
rect -2164 1736 -1964 1783
rect -1906 1817 -1706 1833
rect -1906 1783 -1890 1817
rect -1722 1783 -1706 1817
rect -1906 1736 -1706 1783
rect -1648 1817 -1448 1833
rect -1648 1783 -1632 1817
rect -1464 1783 -1448 1817
rect -1648 1736 -1448 1783
rect -1390 1817 -1190 1833
rect -1390 1783 -1374 1817
rect -1206 1783 -1190 1817
rect -1390 1736 -1190 1783
rect -1132 1817 -932 1833
rect -1132 1783 -1116 1817
rect -948 1783 -932 1817
rect -1132 1736 -932 1783
rect -874 1817 -674 1833
rect -874 1783 -858 1817
rect -690 1783 -674 1817
rect -874 1736 -674 1783
rect -616 1817 -416 1833
rect -616 1783 -600 1817
rect -432 1783 -416 1817
rect -616 1736 -416 1783
rect -358 1817 -158 1833
rect -358 1783 -342 1817
rect -174 1783 -158 1817
rect -358 1736 -158 1783
rect -100 1817 100 1833
rect -100 1783 -84 1817
rect 84 1783 100 1817
rect -100 1736 100 1783
rect 158 1817 358 1833
rect 158 1783 174 1817
rect 342 1783 358 1817
rect 158 1736 358 1783
rect 416 1817 616 1833
rect 416 1783 432 1817
rect 600 1783 616 1817
rect 416 1736 616 1783
rect 674 1817 874 1833
rect 674 1783 690 1817
rect 858 1783 874 1817
rect 674 1736 874 1783
rect 932 1817 1132 1833
rect 932 1783 948 1817
rect 1116 1783 1132 1817
rect 932 1736 1132 1783
rect 1190 1817 1390 1833
rect 1190 1783 1206 1817
rect 1374 1783 1390 1817
rect 1190 1736 1390 1783
rect 1448 1817 1648 1833
rect 1448 1783 1464 1817
rect 1632 1783 1648 1817
rect 1448 1736 1648 1783
rect 1706 1817 1906 1833
rect 1706 1783 1722 1817
rect 1890 1783 1906 1817
rect 1706 1736 1906 1783
rect 1964 1817 2164 1833
rect 1964 1783 1980 1817
rect 2148 1783 2164 1817
rect 1964 1736 2164 1783
rect 2222 1817 2422 1833
rect 2222 1783 2238 1817
rect 2406 1783 2422 1817
rect 2222 1736 2422 1783
rect 2480 1817 2680 1833
rect 2480 1783 2496 1817
rect 2664 1783 2680 1817
rect 2480 1736 2680 1783
rect 2738 1817 2938 1833
rect 2738 1783 2754 1817
rect 2922 1783 2938 1817
rect 2738 1736 2938 1783
rect -2938 689 -2738 736
rect -2938 655 -2922 689
rect -2754 655 -2738 689
rect -2938 639 -2738 655
rect -2680 689 -2480 736
rect -2680 655 -2664 689
rect -2496 655 -2480 689
rect -2680 639 -2480 655
rect -2422 689 -2222 736
rect -2422 655 -2406 689
rect -2238 655 -2222 689
rect -2422 639 -2222 655
rect -2164 689 -1964 736
rect -2164 655 -2148 689
rect -1980 655 -1964 689
rect -2164 639 -1964 655
rect -1906 689 -1706 736
rect -1906 655 -1890 689
rect -1722 655 -1706 689
rect -1906 639 -1706 655
rect -1648 689 -1448 736
rect -1648 655 -1632 689
rect -1464 655 -1448 689
rect -1648 639 -1448 655
rect -1390 689 -1190 736
rect -1390 655 -1374 689
rect -1206 655 -1190 689
rect -1390 639 -1190 655
rect -1132 689 -932 736
rect -1132 655 -1116 689
rect -948 655 -932 689
rect -1132 639 -932 655
rect -874 689 -674 736
rect -874 655 -858 689
rect -690 655 -674 689
rect -874 639 -674 655
rect -616 689 -416 736
rect -616 655 -600 689
rect -432 655 -416 689
rect -616 639 -416 655
rect -358 689 -158 736
rect -358 655 -342 689
rect -174 655 -158 689
rect -358 639 -158 655
rect -100 689 100 736
rect -100 655 -84 689
rect 84 655 100 689
rect -100 639 100 655
rect 158 689 358 736
rect 158 655 174 689
rect 342 655 358 689
rect 158 639 358 655
rect 416 689 616 736
rect 416 655 432 689
rect 600 655 616 689
rect 416 639 616 655
rect 674 689 874 736
rect 674 655 690 689
rect 858 655 874 689
rect 674 639 874 655
rect 932 689 1132 736
rect 932 655 948 689
rect 1116 655 1132 689
rect 932 639 1132 655
rect 1190 689 1390 736
rect 1190 655 1206 689
rect 1374 655 1390 689
rect 1190 639 1390 655
rect 1448 689 1648 736
rect 1448 655 1464 689
rect 1632 655 1648 689
rect 1448 639 1648 655
rect 1706 689 1906 736
rect 1706 655 1722 689
rect 1890 655 1906 689
rect 1706 639 1906 655
rect 1964 689 2164 736
rect 1964 655 1980 689
rect 2148 655 2164 689
rect 1964 639 2164 655
rect 2222 689 2422 736
rect 2222 655 2238 689
rect 2406 655 2422 689
rect 2222 639 2422 655
rect 2480 689 2680 736
rect 2480 655 2496 689
rect 2664 655 2680 689
rect 2480 639 2680 655
rect 2738 689 2938 736
rect 2738 655 2754 689
rect 2922 655 2938 689
rect 2738 639 2938 655
rect -2938 581 -2738 597
rect -2938 547 -2922 581
rect -2754 547 -2738 581
rect -2938 500 -2738 547
rect -2680 581 -2480 597
rect -2680 547 -2664 581
rect -2496 547 -2480 581
rect -2680 500 -2480 547
rect -2422 581 -2222 597
rect -2422 547 -2406 581
rect -2238 547 -2222 581
rect -2422 500 -2222 547
rect -2164 581 -1964 597
rect -2164 547 -2148 581
rect -1980 547 -1964 581
rect -2164 500 -1964 547
rect -1906 581 -1706 597
rect -1906 547 -1890 581
rect -1722 547 -1706 581
rect -1906 500 -1706 547
rect -1648 581 -1448 597
rect -1648 547 -1632 581
rect -1464 547 -1448 581
rect -1648 500 -1448 547
rect -1390 581 -1190 597
rect -1390 547 -1374 581
rect -1206 547 -1190 581
rect -1390 500 -1190 547
rect -1132 581 -932 597
rect -1132 547 -1116 581
rect -948 547 -932 581
rect -1132 500 -932 547
rect -874 581 -674 597
rect -874 547 -858 581
rect -690 547 -674 581
rect -874 500 -674 547
rect -616 581 -416 597
rect -616 547 -600 581
rect -432 547 -416 581
rect -616 500 -416 547
rect -358 581 -158 597
rect -358 547 -342 581
rect -174 547 -158 581
rect -358 500 -158 547
rect -100 581 100 597
rect -100 547 -84 581
rect 84 547 100 581
rect -100 500 100 547
rect 158 581 358 597
rect 158 547 174 581
rect 342 547 358 581
rect 158 500 358 547
rect 416 581 616 597
rect 416 547 432 581
rect 600 547 616 581
rect 416 500 616 547
rect 674 581 874 597
rect 674 547 690 581
rect 858 547 874 581
rect 674 500 874 547
rect 932 581 1132 597
rect 932 547 948 581
rect 1116 547 1132 581
rect 932 500 1132 547
rect 1190 581 1390 597
rect 1190 547 1206 581
rect 1374 547 1390 581
rect 1190 500 1390 547
rect 1448 581 1648 597
rect 1448 547 1464 581
rect 1632 547 1648 581
rect 1448 500 1648 547
rect 1706 581 1906 597
rect 1706 547 1722 581
rect 1890 547 1906 581
rect 1706 500 1906 547
rect 1964 581 2164 597
rect 1964 547 1980 581
rect 2148 547 2164 581
rect 1964 500 2164 547
rect 2222 581 2422 597
rect 2222 547 2238 581
rect 2406 547 2422 581
rect 2222 500 2422 547
rect 2480 581 2680 597
rect 2480 547 2496 581
rect 2664 547 2680 581
rect 2480 500 2680 547
rect 2738 581 2938 597
rect 2738 547 2754 581
rect 2922 547 2938 581
rect 2738 500 2938 547
rect -2938 -547 -2738 -500
rect -2938 -581 -2922 -547
rect -2754 -581 -2738 -547
rect -2938 -597 -2738 -581
rect -2680 -547 -2480 -500
rect -2680 -581 -2664 -547
rect -2496 -581 -2480 -547
rect -2680 -597 -2480 -581
rect -2422 -547 -2222 -500
rect -2422 -581 -2406 -547
rect -2238 -581 -2222 -547
rect -2422 -597 -2222 -581
rect -2164 -547 -1964 -500
rect -2164 -581 -2148 -547
rect -1980 -581 -1964 -547
rect -2164 -597 -1964 -581
rect -1906 -547 -1706 -500
rect -1906 -581 -1890 -547
rect -1722 -581 -1706 -547
rect -1906 -597 -1706 -581
rect -1648 -547 -1448 -500
rect -1648 -581 -1632 -547
rect -1464 -581 -1448 -547
rect -1648 -597 -1448 -581
rect -1390 -547 -1190 -500
rect -1390 -581 -1374 -547
rect -1206 -581 -1190 -547
rect -1390 -597 -1190 -581
rect -1132 -547 -932 -500
rect -1132 -581 -1116 -547
rect -948 -581 -932 -547
rect -1132 -597 -932 -581
rect -874 -547 -674 -500
rect -874 -581 -858 -547
rect -690 -581 -674 -547
rect -874 -597 -674 -581
rect -616 -547 -416 -500
rect -616 -581 -600 -547
rect -432 -581 -416 -547
rect -616 -597 -416 -581
rect -358 -547 -158 -500
rect -358 -581 -342 -547
rect -174 -581 -158 -547
rect -358 -597 -158 -581
rect -100 -547 100 -500
rect -100 -581 -84 -547
rect 84 -581 100 -547
rect -100 -597 100 -581
rect 158 -547 358 -500
rect 158 -581 174 -547
rect 342 -581 358 -547
rect 158 -597 358 -581
rect 416 -547 616 -500
rect 416 -581 432 -547
rect 600 -581 616 -547
rect 416 -597 616 -581
rect 674 -547 874 -500
rect 674 -581 690 -547
rect 858 -581 874 -547
rect 674 -597 874 -581
rect 932 -547 1132 -500
rect 932 -581 948 -547
rect 1116 -581 1132 -547
rect 932 -597 1132 -581
rect 1190 -547 1390 -500
rect 1190 -581 1206 -547
rect 1374 -581 1390 -547
rect 1190 -597 1390 -581
rect 1448 -547 1648 -500
rect 1448 -581 1464 -547
rect 1632 -581 1648 -547
rect 1448 -597 1648 -581
rect 1706 -547 1906 -500
rect 1706 -581 1722 -547
rect 1890 -581 1906 -547
rect 1706 -597 1906 -581
rect 1964 -547 2164 -500
rect 1964 -581 1980 -547
rect 2148 -581 2164 -547
rect 1964 -597 2164 -581
rect 2222 -547 2422 -500
rect 2222 -581 2238 -547
rect 2406 -581 2422 -547
rect 2222 -597 2422 -581
rect 2480 -547 2680 -500
rect 2480 -581 2496 -547
rect 2664 -581 2680 -547
rect 2480 -597 2680 -581
rect 2738 -547 2938 -500
rect 2738 -581 2754 -547
rect 2922 -581 2938 -547
rect 2738 -597 2938 -581
rect -2938 -655 -2738 -639
rect -2938 -689 -2922 -655
rect -2754 -689 -2738 -655
rect -2938 -736 -2738 -689
rect -2680 -655 -2480 -639
rect -2680 -689 -2664 -655
rect -2496 -689 -2480 -655
rect -2680 -736 -2480 -689
rect -2422 -655 -2222 -639
rect -2422 -689 -2406 -655
rect -2238 -689 -2222 -655
rect -2422 -736 -2222 -689
rect -2164 -655 -1964 -639
rect -2164 -689 -2148 -655
rect -1980 -689 -1964 -655
rect -2164 -736 -1964 -689
rect -1906 -655 -1706 -639
rect -1906 -689 -1890 -655
rect -1722 -689 -1706 -655
rect -1906 -736 -1706 -689
rect -1648 -655 -1448 -639
rect -1648 -689 -1632 -655
rect -1464 -689 -1448 -655
rect -1648 -736 -1448 -689
rect -1390 -655 -1190 -639
rect -1390 -689 -1374 -655
rect -1206 -689 -1190 -655
rect -1390 -736 -1190 -689
rect -1132 -655 -932 -639
rect -1132 -689 -1116 -655
rect -948 -689 -932 -655
rect -1132 -736 -932 -689
rect -874 -655 -674 -639
rect -874 -689 -858 -655
rect -690 -689 -674 -655
rect -874 -736 -674 -689
rect -616 -655 -416 -639
rect -616 -689 -600 -655
rect -432 -689 -416 -655
rect -616 -736 -416 -689
rect -358 -655 -158 -639
rect -358 -689 -342 -655
rect -174 -689 -158 -655
rect -358 -736 -158 -689
rect -100 -655 100 -639
rect -100 -689 -84 -655
rect 84 -689 100 -655
rect -100 -736 100 -689
rect 158 -655 358 -639
rect 158 -689 174 -655
rect 342 -689 358 -655
rect 158 -736 358 -689
rect 416 -655 616 -639
rect 416 -689 432 -655
rect 600 -689 616 -655
rect 416 -736 616 -689
rect 674 -655 874 -639
rect 674 -689 690 -655
rect 858 -689 874 -655
rect 674 -736 874 -689
rect 932 -655 1132 -639
rect 932 -689 948 -655
rect 1116 -689 1132 -655
rect 932 -736 1132 -689
rect 1190 -655 1390 -639
rect 1190 -689 1206 -655
rect 1374 -689 1390 -655
rect 1190 -736 1390 -689
rect 1448 -655 1648 -639
rect 1448 -689 1464 -655
rect 1632 -689 1648 -655
rect 1448 -736 1648 -689
rect 1706 -655 1906 -639
rect 1706 -689 1722 -655
rect 1890 -689 1906 -655
rect 1706 -736 1906 -689
rect 1964 -655 2164 -639
rect 1964 -689 1980 -655
rect 2148 -689 2164 -655
rect 1964 -736 2164 -689
rect 2222 -655 2422 -639
rect 2222 -689 2238 -655
rect 2406 -689 2422 -655
rect 2222 -736 2422 -689
rect 2480 -655 2680 -639
rect 2480 -689 2496 -655
rect 2664 -689 2680 -655
rect 2480 -736 2680 -689
rect 2738 -655 2938 -639
rect 2738 -689 2754 -655
rect 2922 -689 2938 -655
rect 2738 -736 2938 -689
rect -2938 -1783 -2738 -1736
rect -2938 -1817 -2922 -1783
rect -2754 -1817 -2738 -1783
rect -2938 -1833 -2738 -1817
rect -2680 -1783 -2480 -1736
rect -2680 -1817 -2664 -1783
rect -2496 -1817 -2480 -1783
rect -2680 -1833 -2480 -1817
rect -2422 -1783 -2222 -1736
rect -2422 -1817 -2406 -1783
rect -2238 -1817 -2222 -1783
rect -2422 -1833 -2222 -1817
rect -2164 -1783 -1964 -1736
rect -2164 -1817 -2148 -1783
rect -1980 -1817 -1964 -1783
rect -2164 -1833 -1964 -1817
rect -1906 -1783 -1706 -1736
rect -1906 -1817 -1890 -1783
rect -1722 -1817 -1706 -1783
rect -1906 -1833 -1706 -1817
rect -1648 -1783 -1448 -1736
rect -1648 -1817 -1632 -1783
rect -1464 -1817 -1448 -1783
rect -1648 -1833 -1448 -1817
rect -1390 -1783 -1190 -1736
rect -1390 -1817 -1374 -1783
rect -1206 -1817 -1190 -1783
rect -1390 -1833 -1190 -1817
rect -1132 -1783 -932 -1736
rect -1132 -1817 -1116 -1783
rect -948 -1817 -932 -1783
rect -1132 -1833 -932 -1817
rect -874 -1783 -674 -1736
rect -874 -1817 -858 -1783
rect -690 -1817 -674 -1783
rect -874 -1833 -674 -1817
rect -616 -1783 -416 -1736
rect -616 -1817 -600 -1783
rect -432 -1817 -416 -1783
rect -616 -1833 -416 -1817
rect -358 -1783 -158 -1736
rect -358 -1817 -342 -1783
rect -174 -1817 -158 -1783
rect -358 -1833 -158 -1817
rect -100 -1783 100 -1736
rect -100 -1817 -84 -1783
rect 84 -1817 100 -1783
rect -100 -1833 100 -1817
rect 158 -1783 358 -1736
rect 158 -1817 174 -1783
rect 342 -1817 358 -1783
rect 158 -1833 358 -1817
rect 416 -1783 616 -1736
rect 416 -1817 432 -1783
rect 600 -1817 616 -1783
rect 416 -1833 616 -1817
rect 674 -1783 874 -1736
rect 674 -1817 690 -1783
rect 858 -1817 874 -1783
rect 674 -1833 874 -1817
rect 932 -1783 1132 -1736
rect 932 -1817 948 -1783
rect 1116 -1817 1132 -1783
rect 932 -1833 1132 -1817
rect 1190 -1783 1390 -1736
rect 1190 -1817 1206 -1783
rect 1374 -1817 1390 -1783
rect 1190 -1833 1390 -1817
rect 1448 -1783 1648 -1736
rect 1448 -1817 1464 -1783
rect 1632 -1817 1648 -1783
rect 1448 -1833 1648 -1817
rect 1706 -1783 1906 -1736
rect 1706 -1817 1722 -1783
rect 1890 -1817 1906 -1783
rect 1706 -1833 1906 -1817
rect 1964 -1783 2164 -1736
rect 1964 -1817 1980 -1783
rect 2148 -1817 2164 -1783
rect 1964 -1833 2164 -1817
rect 2222 -1783 2422 -1736
rect 2222 -1817 2238 -1783
rect 2406 -1817 2422 -1783
rect 2222 -1833 2422 -1817
rect 2480 -1783 2680 -1736
rect 2480 -1817 2496 -1783
rect 2664 -1817 2680 -1783
rect 2480 -1833 2680 -1817
rect 2738 -1783 2938 -1736
rect 2738 -1817 2754 -1783
rect 2922 -1817 2938 -1783
rect 2738 -1833 2938 -1817
rect -2938 -1891 -2738 -1875
rect -2938 -1925 -2922 -1891
rect -2754 -1925 -2738 -1891
rect -2938 -1972 -2738 -1925
rect -2680 -1891 -2480 -1875
rect -2680 -1925 -2664 -1891
rect -2496 -1925 -2480 -1891
rect -2680 -1972 -2480 -1925
rect -2422 -1891 -2222 -1875
rect -2422 -1925 -2406 -1891
rect -2238 -1925 -2222 -1891
rect -2422 -1972 -2222 -1925
rect -2164 -1891 -1964 -1875
rect -2164 -1925 -2148 -1891
rect -1980 -1925 -1964 -1891
rect -2164 -1972 -1964 -1925
rect -1906 -1891 -1706 -1875
rect -1906 -1925 -1890 -1891
rect -1722 -1925 -1706 -1891
rect -1906 -1972 -1706 -1925
rect -1648 -1891 -1448 -1875
rect -1648 -1925 -1632 -1891
rect -1464 -1925 -1448 -1891
rect -1648 -1972 -1448 -1925
rect -1390 -1891 -1190 -1875
rect -1390 -1925 -1374 -1891
rect -1206 -1925 -1190 -1891
rect -1390 -1972 -1190 -1925
rect -1132 -1891 -932 -1875
rect -1132 -1925 -1116 -1891
rect -948 -1925 -932 -1891
rect -1132 -1972 -932 -1925
rect -874 -1891 -674 -1875
rect -874 -1925 -858 -1891
rect -690 -1925 -674 -1891
rect -874 -1972 -674 -1925
rect -616 -1891 -416 -1875
rect -616 -1925 -600 -1891
rect -432 -1925 -416 -1891
rect -616 -1972 -416 -1925
rect -358 -1891 -158 -1875
rect -358 -1925 -342 -1891
rect -174 -1925 -158 -1891
rect -358 -1972 -158 -1925
rect -100 -1891 100 -1875
rect -100 -1925 -84 -1891
rect 84 -1925 100 -1891
rect -100 -1972 100 -1925
rect 158 -1891 358 -1875
rect 158 -1925 174 -1891
rect 342 -1925 358 -1891
rect 158 -1972 358 -1925
rect 416 -1891 616 -1875
rect 416 -1925 432 -1891
rect 600 -1925 616 -1891
rect 416 -1972 616 -1925
rect 674 -1891 874 -1875
rect 674 -1925 690 -1891
rect 858 -1925 874 -1891
rect 674 -1972 874 -1925
rect 932 -1891 1132 -1875
rect 932 -1925 948 -1891
rect 1116 -1925 1132 -1891
rect 932 -1972 1132 -1925
rect 1190 -1891 1390 -1875
rect 1190 -1925 1206 -1891
rect 1374 -1925 1390 -1891
rect 1190 -1972 1390 -1925
rect 1448 -1891 1648 -1875
rect 1448 -1925 1464 -1891
rect 1632 -1925 1648 -1891
rect 1448 -1972 1648 -1925
rect 1706 -1891 1906 -1875
rect 1706 -1925 1722 -1891
rect 1890 -1925 1906 -1891
rect 1706 -1972 1906 -1925
rect 1964 -1891 2164 -1875
rect 1964 -1925 1980 -1891
rect 2148 -1925 2164 -1891
rect 1964 -1972 2164 -1925
rect 2222 -1891 2422 -1875
rect 2222 -1925 2238 -1891
rect 2406 -1925 2422 -1891
rect 2222 -1972 2422 -1925
rect 2480 -1891 2680 -1875
rect 2480 -1925 2496 -1891
rect 2664 -1925 2680 -1891
rect 2480 -1972 2680 -1925
rect 2738 -1891 2938 -1875
rect 2738 -1925 2754 -1891
rect 2922 -1925 2938 -1891
rect 2738 -1972 2938 -1925
rect -2938 -3019 -2738 -2972
rect -2938 -3053 -2922 -3019
rect -2754 -3053 -2738 -3019
rect -2938 -3069 -2738 -3053
rect -2680 -3019 -2480 -2972
rect -2680 -3053 -2664 -3019
rect -2496 -3053 -2480 -3019
rect -2680 -3069 -2480 -3053
rect -2422 -3019 -2222 -2972
rect -2422 -3053 -2406 -3019
rect -2238 -3053 -2222 -3019
rect -2422 -3069 -2222 -3053
rect -2164 -3019 -1964 -2972
rect -2164 -3053 -2148 -3019
rect -1980 -3053 -1964 -3019
rect -2164 -3069 -1964 -3053
rect -1906 -3019 -1706 -2972
rect -1906 -3053 -1890 -3019
rect -1722 -3053 -1706 -3019
rect -1906 -3069 -1706 -3053
rect -1648 -3019 -1448 -2972
rect -1648 -3053 -1632 -3019
rect -1464 -3053 -1448 -3019
rect -1648 -3069 -1448 -3053
rect -1390 -3019 -1190 -2972
rect -1390 -3053 -1374 -3019
rect -1206 -3053 -1190 -3019
rect -1390 -3069 -1190 -3053
rect -1132 -3019 -932 -2972
rect -1132 -3053 -1116 -3019
rect -948 -3053 -932 -3019
rect -1132 -3069 -932 -3053
rect -874 -3019 -674 -2972
rect -874 -3053 -858 -3019
rect -690 -3053 -674 -3019
rect -874 -3069 -674 -3053
rect -616 -3019 -416 -2972
rect -616 -3053 -600 -3019
rect -432 -3053 -416 -3019
rect -616 -3069 -416 -3053
rect -358 -3019 -158 -2972
rect -358 -3053 -342 -3019
rect -174 -3053 -158 -3019
rect -358 -3069 -158 -3053
rect -100 -3019 100 -2972
rect -100 -3053 -84 -3019
rect 84 -3053 100 -3019
rect -100 -3069 100 -3053
rect 158 -3019 358 -2972
rect 158 -3053 174 -3019
rect 342 -3053 358 -3019
rect 158 -3069 358 -3053
rect 416 -3019 616 -2972
rect 416 -3053 432 -3019
rect 600 -3053 616 -3019
rect 416 -3069 616 -3053
rect 674 -3019 874 -2972
rect 674 -3053 690 -3019
rect 858 -3053 874 -3019
rect 674 -3069 874 -3053
rect 932 -3019 1132 -2972
rect 932 -3053 948 -3019
rect 1116 -3053 1132 -3019
rect 932 -3069 1132 -3053
rect 1190 -3019 1390 -2972
rect 1190 -3053 1206 -3019
rect 1374 -3053 1390 -3019
rect 1190 -3069 1390 -3053
rect 1448 -3019 1648 -2972
rect 1448 -3053 1464 -3019
rect 1632 -3053 1648 -3019
rect 1448 -3069 1648 -3053
rect 1706 -3019 1906 -2972
rect 1706 -3053 1722 -3019
rect 1890 -3053 1906 -3019
rect 1706 -3069 1906 -3053
rect 1964 -3019 2164 -2972
rect 1964 -3053 1980 -3019
rect 2148 -3053 2164 -3019
rect 1964 -3069 2164 -3053
rect 2222 -3019 2422 -2972
rect 2222 -3053 2238 -3019
rect 2406 -3053 2422 -3019
rect 2222 -3069 2422 -3053
rect 2480 -3019 2680 -2972
rect 2480 -3053 2496 -3019
rect 2664 -3053 2680 -3019
rect 2480 -3069 2680 -3053
rect 2738 -3019 2938 -2972
rect 2738 -3053 2754 -3019
rect 2922 -3053 2938 -3019
rect 2738 -3069 2938 -3053
<< polycont >>
rect -2922 3019 -2754 3053
rect -2664 3019 -2496 3053
rect -2406 3019 -2238 3053
rect -2148 3019 -1980 3053
rect -1890 3019 -1722 3053
rect -1632 3019 -1464 3053
rect -1374 3019 -1206 3053
rect -1116 3019 -948 3053
rect -858 3019 -690 3053
rect -600 3019 -432 3053
rect -342 3019 -174 3053
rect -84 3019 84 3053
rect 174 3019 342 3053
rect 432 3019 600 3053
rect 690 3019 858 3053
rect 948 3019 1116 3053
rect 1206 3019 1374 3053
rect 1464 3019 1632 3053
rect 1722 3019 1890 3053
rect 1980 3019 2148 3053
rect 2238 3019 2406 3053
rect 2496 3019 2664 3053
rect 2754 3019 2922 3053
rect -2922 1891 -2754 1925
rect -2664 1891 -2496 1925
rect -2406 1891 -2238 1925
rect -2148 1891 -1980 1925
rect -1890 1891 -1722 1925
rect -1632 1891 -1464 1925
rect -1374 1891 -1206 1925
rect -1116 1891 -948 1925
rect -858 1891 -690 1925
rect -600 1891 -432 1925
rect -342 1891 -174 1925
rect -84 1891 84 1925
rect 174 1891 342 1925
rect 432 1891 600 1925
rect 690 1891 858 1925
rect 948 1891 1116 1925
rect 1206 1891 1374 1925
rect 1464 1891 1632 1925
rect 1722 1891 1890 1925
rect 1980 1891 2148 1925
rect 2238 1891 2406 1925
rect 2496 1891 2664 1925
rect 2754 1891 2922 1925
rect -2922 1783 -2754 1817
rect -2664 1783 -2496 1817
rect -2406 1783 -2238 1817
rect -2148 1783 -1980 1817
rect -1890 1783 -1722 1817
rect -1632 1783 -1464 1817
rect -1374 1783 -1206 1817
rect -1116 1783 -948 1817
rect -858 1783 -690 1817
rect -600 1783 -432 1817
rect -342 1783 -174 1817
rect -84 1783 84 1817
rect 174 1783 342 1817
rect 432 1783 600 1817
rect 690 1783 858 1817
rect 948 1783 1116 1817
rect 1206 1783 1374 1817
rect 1464 1783 1632 1817
rect 1722 1783 1890 1817
rect 1980 1783 2148 1817
rect 2238 1783 2406 1817
rect 2496 1783 2664 1817
rect 2754 1783 2922 1817
rect -2922 655 -2754 689
rect -2664 655 -2496 689
rect -2406 655 -2238 689
rect -2148 655 -1980 689
rect -1890 655 -1722 689
rect -1632 655 -1464 689
rect -1374 655 -1206 689
rect -1116 655 -948 689
rect -858 655 -690 689
rect -600 655 -432 689
rect -342 655 -174 689
rect -84 655 84 689
rect 174 655 342 689
rect 432 655 600 689
rect 690 655 858 689
rect 948 655 1116 689
rect 1206 655 1374 689
rect 1464 655 1632 689
rect 1722 655 1890 689
rect 1980 655 2148 689
rect 2238 655 2406 689
rect 2496 655 2664 689
rect 2754 655 2922 689
rect -2922 547 -2754 581
rect -2664 547 -2496 581
rect -2406 547 -2238 581
rect -2148 547 -1980 581
rect -1890 547 -1722 581
rect -1632 547 -1464 581
rect -1374 547 -1206 581
rect -1116 547 -948 581
rect -858 547 -690 581
rect -600 547 -432 581
rect -342 547 -174 581
rect -84 547 84 581
rect 174 547 342 581
rect 432 547 600 581
rect 690 547 858 581
rect 948 547 1116 581
rect 1206 547 1374 581
rect 1464 547 1632 581
rect 1722 547 1890 581
rect 1980 547 2148 581
rect 2238 547 2406 581
rect 2496 547 2664 581
rect 2754 547 2922 581
rect -2922 -581 -2754 -547
rect -2664 -581 -2496 -547
rect -2406 -581 -2238 -547
rect -2148 -581 -1980 -547
rect -1890 -581 -1722 -547
rect -1632 -581 -1464 -547
rect -1374 -581 -1206 -547
rect -1116 -581 -948 -547
rect -858 -581 -690 -547
rect -600 -581 -432 -547
rect -342 -581 -174 -547
rect -84 -581 84 -547
rect 174 -581 342 -547
rect 432 -581 600 -547
rect 690 -581 858 -547
rect 948 -581 1116 -547
rect 1206 -581 1374 -547
rect 1464 -581 1632 -547
rect 1722 -581 1890 -547
rect 1980 -581 2148 -547
rect 2238 -581 2406 -547
rect 2496 -581 2664 -547
rect 2754 -581 2922 -547
rect -2922 -689 -2754 -655
rect -2664 -689 -2496 -655
rect -2406 -689 -2238 -655
rect -2148 -689 -1980 -655
rect -1890 -689 -1722 -655
rect -1632 -689 -1464 -655
rect -1374 -689 -1206 -655
rect -1116 -689 -948 -655
rect -858 -689 -690 -655
rect -600 -689 -432 -655
rect -342 -689 -174 -655
rect -84 -689 84 -655
rect 174 -689 342 -655
rect 432 -689 600 -655
rect 690 -689 858 -655
rect 948 -689 1116 -655
rect 1206 -689 1374 -655
rect 1464 -689 1632 -655
rect 1722 -689 1890 -655
rect 1980 -689 2148 -655
rect 2238 -689 2406 -655
rect 2496 -689 2664 -655
rect 2754 -689 2922 -655
rect -2922 -1817 -2754 -1783
rect -2664 -1817 -2496 -1783
rect -2406 -1817 -2238 -1783
rect -2148 -1817 -1980 -1783
rect -1890 -1817 -1722 -1783
rect -1632 -1817 -1464 -1783
rect -1374 -1817 -1206 -1783
rect -1116 -1817 -948 -1783
rect -858 -1817 -690 -1783
rect -600 -1817 -432 -1783
rect -342 -1817 -174 -1783
rect -84 -1817 84 -1783
rect 174 -1817 342 -1783
rect 432 -1817 600 -1783
rect 690 -1817 858 -1783
rect 948 -1817 1116 -1783
rect 1206 -1817 1374 -1783
rect 1464 -1817 1632 -1783
rect 1722 -1817 1890 -1783
rect 1980 -1817 2148 -1783
rect 2238 -1817 2406 -1783
rect 2496 -1817 2664 -1783
rect 2754 -1817 2922 -1783
rect -2922 -1925 -2754 -1891
rect -2664 -1925 -2496 -1891
rect -2406 -1925 -2238 -1891
rect -2148 -1925 -1980 -1891
rect -1890 -1925 -1722 -1891
rect -1632 -1925 -1464 -1891
rect -1374 -1925 -1206 -1891
rect -1116 -1925 -948 -1891
rect -858 -1925 -690 -1891
rect -600 -1925 -432 -1891
rect -342 -1925 -174 -1891
rect -84 -1925 84 -1891
rect 174 -1925 342 -1891
rect 432 -1925 600 -1891
rect 690 -1925 858 -1891
rect 948 -1925 1116 -1891
rect 1206 -1925 1374 -1891
rect 1464 -1925 1632 -1891
rect 1722 -1925 1890 -1891
rect 1980 -1925 2148 -1891
rect 2238 -1925 2406 -1891
rect 2496 -1925 2664 -1891
rect 2754 -1925 2922 -1891
rect -2922 -3053 -2754 -3019
rect -2664 -3053 -2496 -3019
rect -2406 -3053 -2238 -3019
rect -2148 -3053 -1980 -3019
rect -1890 -3053 -1722 -3019
rect -1632 -3053 -1464 -3019
rect -1374 -3053 -1206 -3019
rect -1116 -3053 -948 -3019
rect -858 -3053 -690 -3019
rect -600 -3053 -432 -3019
rect -342 -3053 -174 -3019
rect -84 -3053 84 -3019
rect 174 -3053 342 -3019
rect 432 -3053 600 -3019
rect 690 -3053 858 -3019
rect 948 -3053 1116 -3019
rect 1206 -3053 1374 -3019
rect 1464 -3053 1632 -3019
rect 1722 -3053 1890 -3019
rect 1980 -3053 2148 -3019
rect 2238 -3053 2406 -3019
rect 2496 -3053 2664 -3019
rect 2754 -3053 2922 -3019
<< locali >>
rect -3118 3157 -3022 3191
rect 3022 3157 3118 3191
rect -3118 3095 -3084 3157
rect 3084 3095 3118 3157
rect -2938 3019 -2922 3053
rect -2754 3019 -2738 3053
rect -2680 3019 -2664 3053
rect -2496 3019 -2480 3053
rect -2422 3019 -2406 3053
rect -2238 3019 -2222 3053
rect -2164 3019 -2148 3053
rect -1980 3019 -1964 3053
rect -1906 3019 -1890 3053
rect -1722 3019 -1706 3053
rect -1648 3019 -1632 3053
rect -1464 3019 -1448 3053
rect -1390 3019 -1374 3053
rect -1206 3019 -1190 3053
rect -1132 3019 -1116 3053
rect -948 3019 -932 3053
rect -874 3019 -858 3053
rect -690 3019 -674 3053
rect -616 3019 -600 3053
rect -432 3019 -416 3053
rect -358 3019 -342 3053
rect -174 3019 -158 3053
rect -100 3019 -84 3053
rect 84 3019 100 3053
rect 158 3019 174 3053
rect 342 3019 358 3053
rect 416 3019 432 3053
rect 600 3019 616 3053
rect 674 3019 690 3053
rect 858 3019 874 3053
rect 932 3019 948 3053
rect 1116 3019 1132 3053
rect 1190 3019 1206 3053
rect 1374 3019 1390 3053
rect 1448 3019 1464 3053
rect 1632 3019 1648 3053
rect 1706 3019 1722 3053
rect 1890 3019 1906 3053
rect 1964 3019 1980 3053
rect 2148 3019 2164 3053
rect 2222 3019 2238 3053
rect 2406 3019 2422 3053
rect 2480 3019 2496 3053
rect 2664 3019 2680 3053
rect 2738 3019 2754 3053
rect 2922 3019 2938 3053
rect -2984 2960 -2950 2976
rect -2984 1968 -2950 1984
rect -2726 2960 -2692 2976
rect -2726 1968 -2692 1984
rect -2468 2960 -2434 2976
rect -2468 1968 -2434 1984
rect -2210 2960 -2176 2976
rect -2210 1968 -2176 1984
rect -1952 2960 -1918 2976
rect -1952 1968 -1918 1984
rect -1694 2960 -1660 2976
rect -1694 1968 -1660 1984
rect -1436 2960 -1402 2976
rect -1436 1968 -1402 1984
rect -1178 2960 -1144 2976
rect -1178 1968 -1144 1984
rect -920 2960 -886 2976
rect -920 1968 -886 1984
rect -662 2960 -628 2976
rect -662 1968 -628 1984
rect -404 2960 -370 2976
rect -404 1968 -370 1984
rect -146 2960 -112 2976
rect -146 1968 -112 1984
rect 112 2960 146 2976
rect 112 1968 146 1984
rect 370 2960 404 2976
rect 370 1968 404 1984
rect 628 2960 662 2976
rect 628 1968 662 1984
rect 886 2960 920 2976
rect 886 1968 920 1984
rect 1144 2960 1178 2976
rect 1144 1968 1178 1984
rect 1402 2960 1436 2976
rect 1402 1968 1436 1984
rect 1660 2960 1694 2976
rect 1660 1968 1694 1984
rect 1918 2960 1952 2976
rect 1918 1968 1952 1984
rect 2176 2960 2210 2976
rect 2176 1968 2210 1984
rect 2434 2960 2468 2976
rect 2434 1968 2468 1984
rect 2692 2960 2726 2976
rect 2692 1968 2726 1984
rect 2950 2960 2984 2976
rect 2950 1968 2984 1984
rect -2938 1891 -2922 1925
rect -2754 1891 -2738 1925
rect -2680 1891 -2664 1925
rect -2496 1891 -2480 1925
rect -2422 1891 -2406 1925
rect -2238 1891 -2222 1925
rect -2164 1891 -2148 1925
rect -1980 1891 -1964 1925
rect -1906 1891 -1890 1925
rect -1722 1891 -1706 1925
rect -1648 1891 -1632 1925
rect -1464 1891 -1448 1925
rect -1390 1891 -1374 1925
rect -1206 1891 -1190 1925
rect -1132 1891 -1116 1925
rect -948 1891 -932 1925
rect -874 1891 -858 1925
rect -690 1891 -674 1925
rect -616 1891 -600 1925
rect -432 1891 -416 1925
rect -358 1891 -342 1925
rect -174 1891 -158 1925
rect -100 1891 -84 1925
rect 84 1891 100 1925
rect 158 1891 174 1925
rect 342 1891 358 1925
rect 416 1891 432 1925
rect 600 1891 616 1925
rect 674 1891 690 1925
rect 858 1891 874 1925
rect 932 1891 948 1925
rect 1116 1891 1132 1925
rect 1190 1891 1206 1925
rect 1374 1891 1390 1925
rect 1448 1891 1464 1925
rect 1632 1891 1648 1925
rect 1706 1891 1722 1925
rect 1890 1891 1906 1925
rect 1964 1891 1980 1925
rect 2148 1891 2164 1925
rect 2222 1891 2238 1925
rect 2406 1891 2422 1925
rect 2480 1891 2496 1925
rect 2664 1891 2680 1925
rect 2738 1891 2754 1925
rect 2922 1891 2938 1925
rect -2938 1783 -2922 1817
rect -2754 1783 -2738 1817
rect -2680 1783 -2664 1817
rect -2496 1783 -2480 1817
rect -2422 1783 -2406 1817
rect -2238 1783 -2222 1817
rect -2164 1783 -2148 1817
rect -1980 1783 -1964 1817
rect -1906 1783 -1890 1817
rect -1722 1783 -1706 1817
rect -1648 1783 -1632 1817
rect -1464 1783 -1448 1817
rect -1390 1783 -1374 1817
rect -1206 1783 -1190 1817
rect -1132 1783 -1116 1817
rect -948 1783 -932 1817
rect -874 1783 -858 1817
rect -690 1783 -674 1817
rect -616 1783 -600 1817
rect -432 1783 -416 1817
rect -358 1783 -342 1817
rect -174 1783 -158 1817
rect -100 1783 -84 1817
rect 84 1783 100 1817
rect 158 1783 174 1817
rect 342 1783 358 1817
rect 416 1783 432 1817
rect 600 1783 616 1817
rect 674 1783 690 1817
rect 858 1783 874 1817
rect 932 1783 948 1817
rect 1116 1783 1132 1817
rect 1190 1783 1206 1817
rect 1374 1783 1390 1817
rect 1448 1783 1464 1817
rect 1632 1783 1648 1817
rect 1706 1783 1722 1817
rect 1890 1783 1906 1817
rect 1964 1783 1980 1817
rect 2148 1783 2164 1817
rect 2222 1783 2238 1817
rect 2406 1783 2422 1817
rect 2480 1783 2496 1817
rect 2664 1783 2680 1817
rect 2738 1783 2754 1817
rect 2922 1783 2938 1817
rect -2984 1724 -2950 1740
rect -2984 732 -2950 748
rect -2726 1724 -2692 1740
rect -2726 732 -2692 748
rect -2468 1724 -2434 1740
rect -2468 732 -2434 748
rect -2210 1724 -2176 1740
rect -2210 732 -2176 748
rect -1952 1724 -1918 1740
rect -1952 732 -1918 748
rect -1694 1724 -1660 1740
rect -1694 732 -1660 748
rect -1436 1724 -1402 1740
rect -1436 732 -1402 748
rect -1178 1724 -1144 1740
rect -1178 732 -1144 748
rect -920 1724 -886 1740
rect -920 732 -886 748
rect -662 1724 -628 1740
rect -662 732 -628 748
rect -404 1724 -370 1740
rect -404 732 -370 748
rect -146 1724 -112 1740
rect -146 732 -112 748
rect 112 1724 146 1740
rect 112 732 146 748
rect 370 1724 404 1740
rect 370 732 404 748
rect 628 1724 662 1740
rect 628 732 662 748
rect 886 1724 920 1740
rect 886 732 920 748
rect 1144 1724 1178 1740
rect 1144 732 1178 748
rect 1402 1724 1436 1740
rect 1402 732 1436 748
rect 1660 1724 1694 1740
rect 1660 732 1694 748
rect 1918 1724 1952 1740
rect 1918 732 1952 748
rect 2176 1724 2210 1740
rect 2176 732 2210 748
rect 2434 1724 2468 1740
rect 2434 732 2468 748
rect 2692 1724 2726 1740
rect 2692 732 2726 748
rect 2950 1724 2984 1740
rect 2950 732 2984 748
rect -2938 655 -2922 689
rect -2754 655 -2738 689
rect -2680 655 -2664 689
rect -2496 655 -2480 689
rect -2422 655 -2406 689
rect -2238 655 -2222 689
rect -2164 655 -2148 689
rect -1980 655 -1964 689
rect -1906 655 -1890 689
rect -1722 655 -1706 689
rect -1648 655 -1632 689
rect -1464 655 -1448 689
rect -1390 655 -1374 689
rect -1206 655 -1190 689
rect -1132 655 -1116 689
rect -948 655 -932 689
rect -874 655 -858 689
rect -690 655 -674 689
rect -616 655 -600 689
rect -432 655 -416 689
rect -358 655 -342 689
rect -174 655 -158 689
rect -100 655 -84 689
rect 84 655 100 689
rect 158 655 174 689
rect 342 655 358 689
rect 416 655 432 689
rect 600 655 616 689
rect 674 655 690 689
rect 858 655 874 689
rect 932 655 948 689
rect 1116 655 1132 689
rect 1190 655 1206 689
rect 1374 655 1390 689
rect 1448 655 1464 689
rect 1632 655 1648 689
rect 1706 655 1722 689
rect 1890 655 1906 689
rect 1964 655 1980 689
rect 2148 655 2164 689
rect 2222 655 2238 689
rect 2406 655 2422 689
rect 2480 655 2496 689
rect 2664 655 2680 689
rect 2738 655 2754 689
rect 2922 655 2938 689
rect -2938 547 -2922 581
rect -2754 547 -2738 581
rect -2680 547 -2664 581
rect -2496 547 -2480 581
rect -2422 547 -2406 581
rect -2238 547 -2222 581
rect -2164 547 -2148 581
rect -1980 547 -1964 581
rect -1906 547 -1890 581
rect -1722 547 -1706 581
rect -1648 547 -1632 581
rect -1464 547 -1448 581
rect -1390 547 -1374 581
rect -1206 547 -1190 581
rect -1132 547 -1116 581
rect -948 547 -932 581
rect -874 547 -858 581
rect -690 547 -674 581
rect -616 547 -600 581
rect -432 547 -416 581
rect -358 547 -342 581
rect -174 547 -158 581
rect -100 547 -84 581
rect 84 547 100 581
rect 158 547 174 581
rect 342 547 358 581
rect 416 547 432 581
rect 600 547 616 581
rect 674 547 690 581
rect 858 547 874 581
rect 932 547 948 581
rect 1116 547 1132 581
rect 1190 547 1206 581
rect 1374 547 1390 581
rect 1448 547 1464 581
rect 1632 547 1648 581
rect 1706 547 1722 581
rect 1890 547 1906 581
rect 1964 547 1980 581
rect 2148 547 2164 581
rect 2222 547 2238 581
rect 2406 547 2422 581
rect 2480 547 2496 581
rect 2664 547 2680 581
rect 2738 547 2754 581
rect 2922 547 2938 581
rect -2984 488 -2950 504
rect -2984 -504 -2950 -488
rect -2726 488 -2692 504
rect -2726 -504 -2692 -488
rect -2468 488 -2434 504
rect -2468 -504 -2434 -488
rect -2210 488 -2176 504
rect -2210 -504 -2176 -488
rect -1952 488 -1918 504
rect -1952 -504 -1918 -488
rect -1694 488 -1660 504
rect -1694 -504 -1660 -488
rect -1436 488 -1402 504
rect -1436 -504 -1402 -488
rect -1178 488 -1144 504
rect -1178 -504 -1144 -488
rect -920 488 -886 504
rect -920 -504 -886 -488
rect -662 488 -628 504
rect -662 -504 -628 -488
rect -404 488 -370 504
rect -404 -504 -370 -488
rect -146 488 -112 504
rect -146 -504 -112 -488
rect 112 488 146 504
rect 112 -504 146 -488
rect 370 488 404 504
rect 370 -504 404 -488
rect 628 488 662 504
rect 628 -504 662 -488
rect 886 488 920 504
rect 886 -504 920 -488
rect 1144 488 1178 504
rect 1144 -504 1178 -488
rect 1402 488 1436 504
rect 1402 -504 1436 -488
rect 1660 488 1694 504
rect 1660 -504 1694 -488
rect 1918 488 1952 504
rect 1918 -504 1952 -488
rect 2176 488 2210 504
rect 2176 -504 2210 -488
rect 2434 488 2468 504
rect 2434 -504 2468 -488
rect 2692 488 2726 504
rect 2692 -504 2726 -488
rect 2950 488 2984 504
rect 2950 -504 2984 -488
rect -2938 -581 -2922 -547
rect -2754 -581 -2738 -547
rect -2680 -581 -2664 -547
rect -2496 -581 -2480 -547
rect -2422 -581 -2406 -547
rect -2238 -581 -2222 -547
rect -2164 -581 -2148 -547
rect -1980 -581 -1964 -547
rect -1906 -581 -1890 -547
rect -1722 -581 -1706 -547
rect -1648 -581 -1632 -547
rect -1464 -581 -1448 -547
rect -1390 -581 -1374 -547
rect -1206 -581 -1190 -547
rect -1132 -581 -1116 -547
rect -948 -581 -932 -547
rect -874 -581 -858 -547
rect -690 -581 -674 -547
rect -616 -581 -600 -547
rect -432 -581 -416 -547
rect -358 -581 -342 -547
rect -174 -581 -158 -547
rect -100 -581 -84 -547
rect 84 -581 100 -547
rect 158 -581 174 -547
rect 342 -581 358 -547
rect 416 -581 432 -547
rect 600 -581 616 -547
rect 674 -581 690 -547
rect 858 -581 874 -547
rect 932 -581 948 -547
rect 1116 -581 1132 -547
rect 1190 -581 1206 -547
rect 1374 -581 1390 -547
rect 1448 -581 1464 -547
rect 1632 -581 1648 -547
rect 1706 -581 1722 -547
rect 1890 -581 1906 -547
rect 1964 -581 1980 -547
rect 2148 -581 2164 -547
rect 2222 -581 2238 -547
rect 2406 -581 2422 -547
rect 2480 -581 2496 -547
rect 2664 -581 2680 -547
rect 2738 -581 2754 -547
rect 2922 -581 2938 -547
rect -2938 -689 -2922 -655
rect -2754 -689 -2738 -655
rect -2680 -689 -2664 -655
rect -2496 -689 -2480 -655
rect -2422 -689 -2406 -655
rect -2238 -689 -2222 -655
rect -2164 -689 -2148 -655
rect -1980 -689 -1964 -655
rect -1906 -689 -1890 -655
rect -1722 -689 -1706 -655
rect -1648 -689 -1632 -655
rect -1464 -689 -1448 -655
rect -1390 -689 -1374 -655
rect -1206 -689 -1190 -655
rect -1132 -689 -1116 -655
rect -948 -689 -932 -655
rect -874 -689 -858 -655
rect -690 -689 -674 -655
rect -616 -689 -600 -655
rect -432 -689 -416 -655
rect -358 -689 -342 -655
rect -174 -689 -158 -655
rect -100 -689 -84 -655
rect 84 -689 100 -655
rect 158 -689 174 -655
rect 342 -689 358 -655
rect 416 -689 432 -655
rect 600 -689 616 -655
rect 674 -689 690 -655
rect 858 -689 874 -655
rect 932 -689 948 -655
rect 1116 -689 1132 -655
rect 1190 -689 1206 -655
rect 1374 -689 1390 -655
rect 1448 -689 1464 -655
rect 1632 -689 1648 -655
rect 1706 -689 1722 -655
rect 1890 -689 1906 -655
rect 1964 -689 1980 -655
rect 2148 -689 2164 -655
rect 2222 -689 2238 -655
rect 2406 -689 2422 -655
rect 2480 -689 2496 -655
rect 2664 -689 2680 -655
rect 2738 -689 2754 -655
rect 2922 -689 2938 -655
rect -2984 -748 -2950 -732
rect -2984 -1740 -2950 -1724
rect -2726 -748 -2692 -732
rect -2726 -1740 -2692 -1724
rect -2468 -748 -2434 -732
rect -2468 -1740 -2434 -1724
rect -2210 -748 -2176 -732
rect -2210 -1740 -2176 -1724
rect -1952 -748 -1918 -732
rect -1952 -1740 -1918 -1724
rect -1694 -748 -1660 -732
rect -1694 -1740 -1660 -1724
rect -1436 -748 -1402 -732
rect -1436 -1740 -1402 -1724
rect -1178 -748 -1144 -732
rect -1178 -1740 -1144 -1724
rect -920 -748 -886 -732
rect -920 -1740 -886 -1724
rect -662 -748 -628 -732
rect -662 -1740 -628 -1724
rect -404 -748 -370 -732
rect -404 -1740 -370 -1724
rect -146 -748 -112 -732
rect -146 -1740 -112 -1724
rect 112 -748 146 -732
rect 112 -1740 146 -1724
rect 370 -748 404 -732
rect 370 -1740 404 -1724
rect 628 -748 662 -732
rect 628 -1740 662 -1724
rect 886 -748 920 -732
rect 886 -1740 920 -1724
rect 1144 -748 1178 -732
rect 1144 -1740 1178 -1724
rect 1402 -748 1436 -732
rect 1402 -1740 1436 -1724
rect 1660 -748 1694 -732
rect 1660 -1740 1694 -1724
rect 1918 -748 1952 -732
rect 1918 -1740 1952 -1724
rect 2176 -748 2210 -732
rect 2176 -1740 2210 -1724
rect 2434 -748 2468 -732
rect 2434 -1740 2468 -1724
rect 2692 -748 2726 -732
rect 2692 -1740 2726 -1724
rect 2950 -748 2984 -732
rect 2950 -1740 2984 -1724
rect -2938 -1817 -2922 -1783
rect -2754 -1817 -2738 -1783
rect -2680 -1817 -2664 -1783
rect -2496 -1817 -2480 -1783
rect -2422 -1817 -2406 -1783
rect -2238 -1817 -2222 -1783
rect -2164 -1817 -2148 -1783
rect -1980 -1817 -1964 -1783
rect -1906 -1817 -1890 -1783
rect -1722 -1817 -1706 -1783
rect -1648 -1817 -1632 -1783
rect -1464 -1817 -1448 -1783
rect -1390 -1817 -1374 -1783
rect -1206 -1817 -1190 -1783
rect -1132 -1817 -1116 -1783
rect -948 -1817 -932 -1783
rect -874 -1817 -858 -1783
rect -690 -1817 -674 -1783
rect -616 -1817 -600 -1783
rect -432 -1817 -416 -1783
rect -358 -1817 -342 -1783
rect -174 -1817 -158 -1783
rect -100 -1817 -84 -1783
rect 84 -1817 100 -1783
rect 158 -1817 174 -1783
rect 342 -1817 358 -1783
rect 416 -1817 432 -1783
rect 600 -1817 616 -1783
rect 674 -1817 690 -1783
rect 858 -1817 874 -1783
rect 932 -1817 948 -1783
rect 1116 -1817 1132 -1783
rect 1190 -1817 1206 -1783
rect 1374 -1817 1390 -1783
rect 1448 -1817 1464 -1783
rect 1632 -1817 1648 -1783
rect 1706 -1817 1722 -1783
rect 1890 -1817 1906 -1783
rect 1964 -1817 1980 -1783
rect 2148 -1817 2164 -1783
rect 2222 -1817 2238 -1783
rect 2406 -1817 2422 -1783
rect 2480 -1817 2496 -1783
rect 2664 -1817 2680 -1783
rect 2738 -1817 2754 -1783
rect 2922 -1817 2938 -1783
rect -2938 -1925 -2922 -1891
rect -2754 -1925 -2738 -1891
rect -2680 -1925 -2664 -1891
rect -2496 -1925 -2480 -1891
rect -2422 -1925 -2406 -1891
rect -2238 -1925 -2222 -1891
rect -2164 -1925 -2148 -1891
rect -1980 -1925 -1964 -1891
rect -1906 -1925 -1890 -1891
rect -1722 -1925 -1706 -1891
rect -1648 -1925 -1632 -1891
rect -1464 -1925 -1448 -1891
rect -1390 -1925 -1374 -1891
rect -1206 -1925 -1190 -1891
rect -1132 -1925 -1116 -1891
rect -948 -1925 -932 -1891
rect -874 -1925 -858 -1891
rect -690 -1925 -674 -1891
rect -616 -1925 -600 -1891
rect -432 -1925 -416 -1891
rect -358 -1925 -342 -1891
rect -174 -1925 -158 -1891
rect -100 -1925 -84 -1891
rect 84 -1925 100 -1891
rect 158 -1925 174 -1891
rect 342 -1925 358 -1891
rect 416 -1925 432 -1891
rect 600 -1925 616 -1891
rect 674 -1925 690 -1891
rect 858 -1925 874 -1891
rect 932 -1925 948 -1891
rect 1116 -1925 1132 -1891
rect 1190 -1925 1206 -1891
rect 1374 -1925 1390 -1891
rect 1448 -1925 1464 -1891
rect 1632 -1925 1648 -1891
rect 1706 -1925 1722 -1891
rect 1890 -1925 1906 -1891
rect 1964 -1925 1980 -1891
rect 2148 -1925 2164 -1891
rect 2222 -1925 2238 -1891
rect 2406 -1925 2422 -1891
rect 2480 -1925 2496 -1891
rect 2664 -1925 2680 -1891
rect 2738 -1925 2754 -1891
rect 2922 -1925 2938 -1891
rect -2984 -1984 -2950 -1968
rect -2984 -2976 -2950 -2960
rect -2726 -1984 -2692 -1968
rect -2726 -2976 -2692 -2960
rect -2468 -1984 -2434 -1968
rect -2468 -2976 -2434 -2960
rect -2210 -1984 -2176 -1968
rect -2210 -2976 -2176 -2960
rect -1952 -1984 -1918 -1968
rect -1952 -2976 -1918 -2960
rect -1694 -1984 -1660 -1968
rect -1694 -2976 -1660 -2960
rect -1436 -1984 -1402 -1968
rect -1436 -2976 -1402 -2960
rect -1178 -1984 -1144 -1968
rect -1178 -2976 -1144 -2960
rect -920 -1984 -886 -1968
rect -920 -2976 -886 -2960
rect -662 -1984 -628 -1968
rect -662 -2976 -628 -2960
rect -404 -1984 -370 -1968
rect -404 -2976 -370 -2960
rect -146 -1984 -112 -1968
rect -146 -2976 -112 -2960
rect 112 -1984 146 -1968
rect 112 -2976 146 -2960
rect 370 -1984 404 -1968
rect 370 -2976 404 -2960
rect 628 -1984 662 -1968
rect 628 -2976 662 -2960
rect 886 -1984 920 -1968
rect 886 -2976 920 -2960
rect 1144 -1984 1178 -1968
rect 1144 -2976 1178 -2960
rect 1402 -1984 1436 -1968
rect 1402 -2976 1436 -2960
rect 1660 -1984 1694 -1968
rect 1660 -2976 1694 -2960
rect 1918 -1984 1952 -1968
rect 1918 -2976 1952 -2960
rect 2176 -1984 2210 -1968
rect 2176 -2976 2210 -2960
rect 2434 -1984 2468 -1968
rect 2434 -2976 2468 -2960
rect 2692 -1984 2726 -1968
rect 2692 -2976 2726 -2960
rect 2950 -1984 2984 -1968
rect 2950 -2976 2984 -2960
rect -2938 -3053 -2922 -3019
rect -2754 -3053 -2738 -3019
rect -2680 -3053 -2664 -3019
rect -2496 -3053 -2480 -3019
rect -2422 -3053 -2406 -3019
rect -2238 -3053 -2222 -3019
rect -2164 -3053 -2148 -3019
rect -1980 -3053 -1964 -3019
rect -1906 -3053 -1890 -3019
rect -1722 -3053 -1706 -3019
rect -1648 -3053 -1632 -3019
rect -1464 -3053 -1448 -3019
rect -1390 -3053 -1374 -3019
rect -1206 -3053 -1190 -3019
rect -1132 -3053 -1116 -3019
rect -948 -3053 -932 -3019
rect -874 -3053 -858 -3019
rect -690 -3053 -674 -3019
rect -616 -3053 -600 -3019
rect -432 -3053 -416 -3019
rect -358 -3053 -342 -3019
rect -174 -3053 -158 -3019
rect -100 -3053 -84 -3019
rect 84 -3053 100 -3019
rect 158 -3053 174 -3019
rect 342 -3053 358 -3019
rect 416 -3053 432 -3019
rect 600 -3053 616 -3019
rect 674 -3053 690 -3019
rect 858 -3053 874 -3019
rect 932 -3053 948 -3019
rect 1116 -3053 1132 -3019
rect 1190 -3053 1206 -3019
rect 1374 -3053 1390 -3019
rect 1448 -3053 1464 -3019
rect 1632 -3053 1648 -3019
rect 1706 -3053 1722 -3019
rect 1890 -3053 1906 -3019
rect 1964 -3053 1980 -3019
rect 2148 -3053 2164 -3019
rect 2222 -3053 2238 -3019
rect 2406 -3053 2422 -3019
rect 2480 -3053 2496 -3019
rect 2664 -3053 2680 -3019
rect 2738 -3053 2754 -3019
rect 2922 -3053 2938 -3019
rect -3118 -3157 -3084 -3095
rect 3084 -3157 3118 -3095
rect -3118 -3191 -3022 -3157
rect 3022 -3191 3118 -3157
<< viali >>
rect -2922 3019 -2754 3053
rect -2664 3019 -2496 3053
rect -2406 3019 -2238 3053
rect -2148 3019 -1980 3053
rect -1890 3019 -1722 3053
rect -1632 3019 -1464 3053
rect -1374 3019 -1206 3053
rect -1116 3019 -948 3053
rect -858 3019 -690 3053
rect -600 3019 -432 3053
rect -342 3019 -174 3053
rect -84 3019 84 3053
rect 174 3019 342 3053
rect 432 3019 600 3053
rect 690 3019 858 3053
rect 948 3019 1116 3053
rect 1206 3019 1374 3053
rect 1464 3019 1632 3053
rect 1722 3019 1890 3053
rect 1980 3019 2148 3053
rect 2238 3019 2406 3053
rect 2496 3019 2664 3053
rect 2754 3019 2922 3053
rect -2984 1984 -2950 2960
rect -2726 1984 -2692 2960
rect -2468 1984 -2434 2960
rect -2210 1984 -2176 2960
rect -1952 1984 -1918 2960
rect -1694 1984 -1660 2960
rect -1436 1984 -1402 2960
rect -1178 1984 -1144 2960
rect -920 1984 -886 2960
rect -662 1984 -628 2960
rect -404 1984 -370 2960
rect -146 1984 -112 2960
rect 112 1984 146 2960
rect 370 1984 404 2960
rect 628 1984 662 2960
rect 886 1984 920 2960
rect 1144 1984 1178 2960
rect 1402 1984 1436 2960
rect 1660 1984 1694 2960
rect 1918 1984 1952 2960
rect 2176 1984 2210 2960
rect 2434 1984 2468 2960
rect 2692 1984 2726 2960
rect 2950 1984 2984 2960
rect -2922 1891 -2754 1925
rect -2664 1891 -2496 1925
rect -2406 1891 -2238 1925
rect -2148 1891 -1980 1925
rect -1890 1891 -1722 1925
rect -1632 1891 -1464 1925
rect -1374 1891 -1206 1925
rect -1116 1891 -948 1925
rect -858 1891 -690 1925
rect -600 1891 -432 1925
rect -342 1891 -174 1925
rect -84 1891 84 1925
rect 174 1891 342 1925
rect 432 1891 600 1925
rect 690 1891 858 1925
rect 948 1891 1116 1925
rect 1206 1891 1374 1925
rect 1464 1891 1632 1925
rect 1722 1891 1890 1925
rect 1980 1891 2148 1925
rect 2238 1891 2406 1925
rect 2496 1891 2664 1925
rect 2754 1891 2922 1925
rect -2922 1783 -2754 1817
rect -2664 1783 -2496 1817
rect -2406 1783 -2238 1817
rect -2148 1783 -1980 1817
rect -1890 1783 -1722 1817
rect -1632 1783 -1464 1817
rect -1374 1783 -1206 1817
rect -1116 1783 -948 1817
rect -858 1783 -690 1817
rect -600 1783 -432 1817
rect -342 1783 -174 1817
rect -84 1783 84 1817
rect 174 1783 342 1817
rect 432 1783 600 1817
rect 690 1783 858 1817
rect 948 1783 1116 1817
rect 1206 1783 1374 1817
rect 1464 1783 1632 1817
rect 1722 1783 1890 1817
rect 1980 1783 2148 1817
rect 2238 1783 2406 1817
rect 2496 1783 2664 1817
rect 2754 1783 2922 1817
rect -2984 748 -2950 1724
rect -2726 748 -2692 1724
rect -2468 748 -2434 1724
rect -2210 748 -2176 1724
rect -1952 748 -1918 1724
rect -1694 748 -1660 1724
rect -1436 748 -1402 1724
rect -1178 748 -1144 1724
rect -920 748 -886 1724
rect -662 748 -628 1724
rect -404 748 -370 1724
rect -146 748 -112 1724
rect 112 748 146 1724
rect 370 748 404 1724
rect 628 748 662 1724
rect 886 748 920 1724
rect 1144 748 1178 1724
rect 1402 748 1436 1724
rect 1660 748 1694 1724
rect 1918 748 1952 1724
rect 2176 748 2210 1724
rect 2434 748 2468 1724
rect 2692 748 2726 1724
rect 2950 748 2984 1724
rect -2922 655 -2754 689
rect -2664 655 -2496 689
rect -2406 655 -2238 689
rect -2148 655 -1980 689
rect -1890 655 -1722 689
rect -1632 655 -1464 689
rect -1374 655 -1206 689
rect -1116 655 -948 689
rect -858 655 -690 689
rect -600 655 -432 689
rect -342 655 -174 689
rect -84 655 84 689
rect 174 655 342 689
rect 432 655 600 689
rect 690 655 858 689
rect 948 655 1116 689
rect 1206 655 1374 689
rect 1464 655 1632 689
rect 1722 655 1890 689
rect 1980 655 2148 689
rect 2238 655 2406 689
rect 2496 655 2664 689
rect 2754 655 2922 689
rect -2922 547 -2754 581
rect -2664 547 -2496 581
rect -2406 547 -2238 581
rect -2148 547 -1980 581
rect -1890 547 -1722 581
rect -1632 547 -1464 581
rect -1374 547 -1206 581
rect -1116 547 -948 581
rect -858 547 -690 581
rect -600 547 -432 581
rect -342 547 -174 581
rect -84 547 84 581
rect 174 547 342 581
rect 432 547 600 581
rect 690 547 858 581
rect 948 547 1116 581
rect 1206 547 1374 581
rect 1464 547 1632 581
rect 1722 547 1890 581
rect 1980 547 2148 581
rect 2238 547 2406 581
rect 2496 547 2664 581
rect 2754 547 2922 581
rect -2984 -488 -2950 488
rect -2726 -488 -2692 488
rect -2468 -488 -2434 488
rect -2210 -488 -2176 488
rect -1952 -488 -1918 488
rect -1694 -488 -1660 488
rect -1436 -488 -1402 488
rect -1178 -488 -1144 488
rect -920 -488 -886 488
rect -662 -488 -628 488
rect -404 -488 -370 488
rect -146 -488 -112 488
rect 112 -488 146 488
rect 370 -488 404 488
rect 628 -488 662 488
rect 886 -488 920 488
rect 1144 -488 1178 488
rect 1402 -488 1436 488
rect 1660 -488 1694 488
rect 1918 -488 1952 488
rect 2176 -488 2210 488
rect 2434 -488 2468 488
rect 2692 -488 2726 488
rect 2950 -488 2984 488
rect -2922 -581 -2754 -547
rect -2664 -581 -2496 -547
rect -2406 -581 -2238 -547
rect -2148 -581 -1980 -547
rect -1890 -581 -1722 -547
rect -1632 -581 -1464 -547
rect -1374 -581 -1206 -547
rect -1116 -581 -948 -547
rect -858 -581 -690 -547
rect -600 -581 -432 -547
rect -342 -581 -174 -547
rect -84 -581 84 -547
rect 174 -581 342 -547
rect 432 -581 600 -547
rect 690 -581 858 -547
rect 948 -581 1116 -547
rect 1206 -581 1374 -547
rect 1464 -581 1632 -547
rect 1722 -581 1890 -547
rect 1980 -581 2148 -547
rect 2238 -581 2406 -547
rect 2496 -581 2664 -547
rect 2754 -581 2922 -547
rect -2922 -689 -2754 -655
rect -2664 -689 -2496 -655
rect -2406 -689 -2238 -655
rect -2148 -689 -1980 -655
rect -1890 -689 -1722 -655
rect -1632 -689 -1464 -655
rect -1374 -689 -1206 -655
rect -1116 -689 -948 -655
rect -858 -689 -690 -655
rect -600 -689 -432 -655
rect -342 -689 -174 -655
rect -84 -689 84 -655
rect 174 -689 342 -655
rect 432 -689 600 -655
rect 690 -689 858 -655
rect 948 -689 1116 -655
rect 1206 -689 1374 -655
rect 1464 -689 1632 -655
rect 1722 -689 1890 -655
rect 1980 -689 2148 -655
rect 2238 -689 2406 -655
rect 2496 -689 2664 -655
rect 2754 -689 2922 -655
rect -2984 -1724 -2950 -748
rect -2726 -1724 -2692 -748
rect -2468 -1724 -2434 -748
rect -2210 -1724 -2176 -748
rect -1952 -1724 -1918 -748
rect -1694 -1724 -1660 -748
rect -1436 -1724 -1402 -748
rect -1178 -1724 -1144 -748
rect -920 -1724 -886 -748
rect -662 -1724 -628 -748
rect -404 -1724 -370 -748
rect -146 -1724 -112 -748
rect 112 -1724 146 -748
rect 370 -1724 404 -748
rect 628 -1724 662 -748
rect 886 -1724 920 -748
rect 1144 -1724 1178 -748
rect 1402 -1724 1436 -748
rect 1660 -1724 1694 -748
rect 1918 -1724 1952 -748
rect 2176 -1724 2210 -748
rect 2434 -1724 2468 -748
rect 2692 -1724 2726 -748
rect 2950 -1724 2984 -748
rect -2922 -1817 -2754 -1783
rect -2664 -1817 -2496 -1783
rect -2406 -1817 -2238 -1783
rect -2148 -1817 -1980 -1783
rect -1890 -1817 -1722 -1783
rect -1632 -1817 -1464 -1783
rect -1374 -1817 -1206 -1783
rect -1116 -1817 -948 -1783
rect -858 -1817 -690 -1783
rect -600 -1817 -432 -1783
rect -342 -1817 -174 -1783
rect -84 -1817 84 -1783
rect 174 -1817 342 -1783
rect 432 -1817 600 -1783
rect 690 -1817 858 -1783
rect 948 -1817 1116 -1783
rect 1206 -1817 1374 -1783
rect 1464 -1817 1632 -1783
rect 1722 -1817 1890 -1783
rect 1980 -1817 2148 -1783
rect 2238 -1817 2406 -1783
rect 2496 -1817 2664 -1783
rect 2754 -1817 2922 -1783
rect -2922 -1925 -2754 -1891
rect -2664 -1925 -2496 -1891
rect -2406 -1925 -2238 -1891
rect -2148 -1925 -1980 -1891
rect -1890 -1925 -1722 -1891
rect -1632 -1925 -1464 -1891
rect -1374 -1925 -1206 -1891
rect -1116 -1925 -948 -1891
rect -858 -1925 -690 -1891
rect -600 -1925 -432 -1891
rect -342 -1925 -174 -1891
rect -84 -1925 84 -1891
rect 174 -1925 342 -1891
rect 432 -1925 600 -1891
rect 690 -1925 858 -1891
rect 948 -1925 1116 -1891
rect 1206 -1925 1374 -1891
rect 1464 -1925 1632 -1891
rect 1722 -1925 1890 -1891
rect 1980 -1925 2148 -1891
rect 2238 -1925 2406 -1891
rect 2496 -1925 2664 -1891
rect 2754 -1925 2922 -1891
rect -2984 -2960 -2950 -1984
rect -2726 -2960 -2692 -1984
rect -2468 -2960 -2434 -1984
rect -2210 -2960 -2176 -1984
rect -1952 -2960 -1918 -1984
rect -1694 -2960 -1660 -1984
rect -1436 -2960 -1402 -1984
rect -1178 -2960 -1144 -1984
rect -920 -2960 -886 -1984
rect -662 -2960 -628 -1984
rect -404 -2960 -370 -1984
rect -146 -2960 -112 -1984
rect 112 -2960 146 -1984
rect 370 -2960 404 -1984
rect 628 -2960 662 -1984
rect 886 -2960 920 -1984
rect 1144 -2960 1178 -1984
rect 1402 -2960 1436 -1984
rect 1660 -2960 1694 -1984
rect 1918 -2960 1952 -1984
rect 2176 -2960 2210 -1984
rect 2434 -2960 2468 -1984
rect 2692 -2960 2726 -1984
rect 2950 -2960 2984 -1984
rect -2922 -3053 -2754 -3019
rect -2664 -3053 -2496 -3019
rect -2406 -3053 -2238 -3019
rect -2148 -3053 -1980 -3019
rect -1890 -3053 -1722 -3019
rect -1632 -3053 -1464 -3019
rect -1374 -3053 -1206 -3019
rect -1116 -3053 -948 -3019
rect -858 -3053 -690 -3019
rect -600 -3053 -432 -3019
rect -342 -3053 -174 -3019
rect -84 -3053 84 -3019
rect 174 -3053 342 -3019
rect 432 -3053 600 -3019
rect 690 -3053 858 -3019
rect 948 -3053 1116 -3019
rect 1206 -3053 1374 -3019
rect 1464 -3053 1632 -3019
rect 1722 -3053 1890 -3019
rect 1980 -3053 2148 -3019
rect 2238 -3053 2406 -3019
rect 2496 -3053 2664 -3019
rect 2754 -3053 2922 -3019
<< metal1 >>
rect -2934 3053 -2742 3059
rect -2934 3019 -2922 3053
rect -2754 3019 -2742 3053
rect -2934 3013 -2742 3019
rect -2676 3053 -2484 3059
rect -2676 3019 -2664 3053
rect -2496 3019 -2484 3053
rect -2676 3013 -2484 3019
rect -2418 3053 -2226 3059
rect -2418 3019 -2406 3053
rect -2238 3019 -2226 3053
rect -2418 3013 -2226 3019
rect -2160 3053 -1968 3059
rect -2160 3019 -2148 3053
rect -1980 3019 -1968 3053
rect -2160 3013 -1968 3019
rect -1902 3053 -1710 3059
rect -1902 3019 -1890 3053
rect -1722 3019 -1710 3053
rect -1902 3013 -1710 3019
rect -1644 3053 -1452 3059
rect -1644 3019 -1632 3053
rect -1464 3019 -1452 3053
rect -1644 3013 -1452 3019
rect -1386 3053 -1194 3059
rect -1386 3019 -1374 3053
rect -1206 3019 -1194 3053
rect -1386 3013 -1194 3019
rect -1128 3053 -936 3059
rect -1128 3019 -1116 3053
rect -948 3019 -936 3053
rect -1128 3013 -936 3019
rect -870 3053 -678 3059
rect -870 3019 -858 3053
rect -690 3019 -678 3053
rect -870 3013 -678 3019
rect -612 3053 -420 3059
rect -612 3019 -600 3053
rect -432 3019 -420 3053
rect -612 3013 -420 3019
rect -354 3053 -162 3059
rect -354 3019 -342 3053
rect -174 3019 -162 3053
rect -354 3013 -162 3019
rect -96 3053 96 3059
rect -96 3019 -84 3053
rect 84 3019 96 3053
rect -96 3013 96 3019
rect 162 3053 354 3059
rect 162 3019 174 3053
rect 342 3019 354 3053
rect 162 3013 354 3019
rect 420 3053 612 3059
rect 420 3019 432 3053
rect 600 3019 612 3053
rect 420 3013 612 3019
rect 678 3053 870 3059
rect 678 3019 690 3053
rect 858 3019 870 3053
rect 678 3013 870 3019
rect 936 3053 1128 3059
rect 936 3019 948 3053
rect 1116 3019 1128 3053
rect 936 3013 1128 3019
rect 1194 3053 1386 3059
rect 1194 3019 1206 3053
rect 1374 3019 1386 3053
rect 1194 3013 1386 3019
rect 1452 3053 1644 3059
rect 1452 3019 1464 3053
rect 1632 3019 1644 3053
rect 1452 3013 1644 3019
rect 1710 3053 1902 3059
rect 1710 3019 1722 3053
rect 1890 3019 1902 3053
rect 1710 3013 1902 3019
rect 1968 3053 2160 3059
rect 1968 3019 1980 3053
rect 2148 3019 2160 3053
rect 1968 3013 2160 3019
rect 2226 3053 2418 3059
rect 2226 3019 2238 3053
rect 2406 3019 2418 3053
rect 2226 3013 2418 3019
rect 2484 3053 2676 3059
rect 2484 3019 2496 3053
rect 2664 3019 2676 3053
rect 2484 3013 2676 3019
rect 2742 3053 2934 3059
rect 2742 3019 2754 3053
rect 2922 3019 2934 3053
rect 2742 3013 2934 3019
rect -2990 2960 -2944 2972
rect -2990 1984 -2984 2960
rect -2950 1984 -2944 2960
rect -2990 1972 -2944 1984
rect -2732 2960 -2686 2972
rect -2732 1984 -2726 2960
rect -2692 1984 -2686 2960
rect -2732 1972 -2686 1984
rect -2474 2960 -2428 2972
rect -2474 1984 -2468 2960
rect -2434 1984 -2428 2960
rect -2474 1972 -2428 1984
rect -2216 2960 -2170 2972
rect -2216 1984 -2210 2960
rect -2176 1984 -2170 2960
rect -2216 1972 -2170 1984
rect -1958 2960 -1912 2972
rect -1958 1984 -1952 2960
rect -1918 1984 -1912 2960
rect -1958 1972 -1912 1984
rect -1700 2960 -1654 2972
rect -1700 1984 -1694 2960
rect -1660 1984 -1654 2960
rect -1700 1972 -1654 1984
rect -1442 2960 -1396 2972
rect -1442 1984 -1436 2960
rect -1402 1984 -1396 2960
rect -1442 1972 -1396 1984
rect -1184 2960 -1138 2972
rect -1184 1984 -1178 2960
rect -1144 1984 -1138 2960
rect -1184 1972 -1138 1984
rect -926 2960 -880 2972
rect -926 1984 -920 2960
rect -886 1984 -880 2960
rect -926 1972 -880 1984
rect -668 2960 -622 2972
rect -668 1984 -662 2960
rect -628 1984 -622 2960
rect -668 1972 -622 1984
rect -410 2960 -364 2972
rect -410 1984 -404 2960
rect -370 1984 -364 2960
rect -410 1972 -364 1984
rect -152 2960 -106 2972
rect -152 1984 -146 2960
rect -112 1984 -106 2960
rect -152 1972 -106 1984
rect 106 2960 152 2972
rect 106 1984 112 2960
rect 146 1984 152 2960
rect 106 1972 152 1984
rect 364 2960 410 2972
rect 364 1984 370 2960
rect 404 1984 410 2960
rect 364 1972 410 1984
rect 622 2960 668 2972
rect 622 1984 628 2960
rect 662 1984 668 2960
rect 622 1972 668 1984
rect 880 2960 926 2972
rect 880 1984 886 2960
rect 920 1984 926 2960
rect 880 1972 926 1984
rect 1138 2960 1184 2972
rect 1138 1984 1144 2960
rect 1178 1984 1184 2960
rect 1138 1972 1184 1984
rect 1396 2960 1442 2972
rect 1396 1984 1402 2960
rect 1436 1984 1442 2960
rect 1396 1972 1442 1984
rect 1654 2960 1700 2972
rect 1654 1984 1660 2960
rect 1694 1984 1700 2960
rect 1654 1972 1700 1984
rect 1912 2960 1958 2972
rect 1912 1984 1918 2960
rect 1952 1984 1958 2960
rect 1912 1972 1958 1984
rect 2170 2960 2216 2972
rect 2170 1984 2176 2960
rect 2210 1984 2216 2960
rect 2170 1972 2216 1984
rect 2428 2960 2474 2972
rect 2428 1984 2434 2960
rect 2468 1984 2474 2960
rect 2428 1972 2474 1984
rect 2686 2960 2732 2972
rect 2686 1984 2692 2960
rect 2726 1984 2732 2960
rect 2686 1972 2732 1984
rect 2944 2960 2990 2972
rect 2944 1984 2950 2960
rect 2984 1984 2990 2960
rect 2944 1972 2990 1984
rect -2934 1925 -2742 1931
rect -2934 1891 -2922 1925
rect -2754 1891 -2742 1925
rect -2934 1885 -2742 1891
rect -2676 1925 -2484 1931
rect -2676 1891 -2664 1925
rect -2496 1891 -2484 1925
rect -2676 1885 -2484 1891
rect -2418 1925 -2226 1931
rect -2418 1891 -2406 1925
rect -2238 1891 -2226 1925
rect -2418 1885 -2226 1891
rect -2160 1925 -1968 1931
rect -2160 1891 -2148 1925
rect -1980 1891 -1968 1925
rect -2160 1885 -1968 1891
rect -1902 1925 -1710 1931
rect -1902 1891 -1890 1925
rect -1722 1891 -1710 1925
rect -1902 1885 -1710 1891
rect -1644 1925 -1452 1931
rect -1644 1891 -1632 1925
rect -1464 1891 -1452 1925
rect -1644 1885 -1452 1891
rect -1386 1925 -1194 1931
rect -1386 1891 -1374 1925
rect -1206 1891 -1194 1925
rect -1386 1885 -1194 1891
rect -1128 1925 -936 1931
rect -1128 1891 -1116 1925
rect -948 1891 -936 1925
rect -1128 1885 -936 1891
rect -870 1925 -678 1931
rect -870 1891 -858 1925
rect -690 1891 -678 1925
rect -870 1885 -678 1891
rect -612 1925 -420 1931
rect -612 1891 -600 1925
rect -432 1891 -420 1925
rect -612 1885 -420 1891
rect -354 1925 -162 1931
rect -354 1891 -342 1925
rect -174 1891 -162 1925
rect -354 1885 -162 1891
rect -96 1925 96 1931
rect -96 1891 -84 1925
rect 84 1891 96 1925
rect -96 1885 96 1891
rect 162 1925 354 1931
rect 162 1891 174 1925
rect 342 1891 354 1925
rect 162 1885 354 1891
rect 420 1925 612 1931
rect 420 1891 432 1925
rect 600 1891 612 1925
rect 420 1885 612 1891
rect 678 1925 870 1931
rect 678 1891 690 1925
rect 858 1891 870 1925
rect 678 1885 870 1891
rect 936 1925 1128 1931
rect 936 1891 948 1925
rect 1116 1891 1128 1925
rect 936 1885 1128 1891
rect 1194 1925 1386 1931
rect 1194 1891 1206 1925
rect 1374 1891 1386 1925
rect 1194 1885 1386 1891
rect 1452 1925 1644 1931
rect 1452 1891 1464 1925
rect 1632 1891 1644 1925
rect 1452 1885 1644 1891
rect 1710 1925 1902 1931
rect 1710 1891 1722 1925
rect 1890 1891 1902 1925
rect 1710 1885 1902 1891
rect 1968 1925 2160 1931
rect 1968 1891 1980 1925
rect 2148 1891 2160 1925
rect 1968 1885 2160 1891
rect 2226 1925 2418 1931
rect 2226 1891 2238 1925
rect 2406 1891 2418 1925
rect 2226 1885 2418 1891
rect 2484 1925 2676 1931
rect 2484 1891 2496 1925
rect 2664 1891 2676 1925
rect 2484 1885 2676 1891
rect 2742 1925 2934 1931
rect 2742 1891 2754 1925
rect 2922 1891 2934 1925
rect 2742 1885 2934 1891
rect -2934 1817 -2742 1823
rect -2934 1783 -2922 1817
rect -2754 1783 -2742 1817
rect -2934 1777 -2742 1783
rect -2676 1817 -2484 1823
rect -2676 1783 -2664 1817
rect -2496 1783 -2484 1817
rect -2676 1777 -2484 1783
rect -2418 1817 -2226 1823
rect -2418 1783 -2406 1817
rect -2238 1783 -2226 1817
rect -2418 1777 -2226 1783
rect -2160 1817 -1968 1823
rect -2160 1783 -2148 1817
rect -1980 1783 -1968 1817
rect -2160 1777 -1968 1783
rect -1902 1817 -1710 1823
rect -1902 1783 -1890 1817
rect -1722 1783 -1710 1817
rect -1902 1777 -1710 1783
rect -1644 1817 -1452 1823
rect -1644 1783 -1632 1817
rect -1464 1783 -1452 1817
rect -1644 1777 -1452 1783
rect -1386 1817 -1194 1823
rect -1386 1783 -1374 1817
rect -1206 1783 -1194 1817
rect -1386 1777 -1194 1783
rect -1128 1817 -936 1823
rect -1128 1783 -1116 1817
rect -948 1783 -936 1817
rect -1128 1777 -936 1783
rect -870 1817 -678 1823
rect -870 1783 -858 1817
rect -690 1783 -678 1817
rect -870 1777 -678 1783
rect -612 1817 -420 1823
rect -612 1783 -600 1817
rect -432 1783 -420 1817
rect -612 1777 -420 1783
rect -354 1817 -162 1823
rect -354 1783 -342 1817
rect -174 1783 -162 1817
rect -354 1777 -162 1783
rect -96 1817 96 1823
rect -96 1783 -84 1817
rect 84 1783 96 1817
rect -96 1777 96 1783
rect 162 1817 354 1823
rect 162 1783 174 1817
rect 342 1783 354 1817
rect 162 1777 354 1783
rect 420 1817 612 1823
rect 420 1783 432 1817
rect 600 1783 612 1817
rect 420 1777 612 1783
rect 678 1817 870 1823
rect 678 1783 690 1817
rect 858 1783 870 1817
rect 678 1777 870 1783
rect 936 1817 1128 1823
rect 936 1783 948 1817
rect 1116 1783 1128 1817
rect 936 1777 1128 1783
rect 1194 1817 1386 1823
rect 1194 1783 1206 1817
rect 1374 1783 1386 1817
rect 1194 1777 1386 1783
rect 1452 1817 1644 1823
rect 1452 1783 1464 1817
rect 1632 1783 1644 1817
rect 1452 1777 1644 1783
rect 1710 1817 1902 1823
rect 1710 1783 1722 1817
rect 1890 1783 1902 1817
rect 1710 1777 1902 1783
rect 1968 1817 2160 1823
rect 1968 1783 1980 1817
rect 2148 1783 2160 1817
rect 1968 1777 2160 1783
rect 2226 1817 2418 1823
rect 2226 1783 2238 1817
rect 2406 1783 2418 1817
rect 2226 1777 2418 1783
rect 2484 1817 2676 1823
rect 2484 1783 2496 1817
rect 2664 1783 2676 1817
rect 2484 1777 2676 1783
rect 2742 1817 2934 1823
rect 2742 1783 2754 1817
rect 2922 1783 2934 1817
rect 2742 1777 2934 1783
rect -2990 1724 -2944 1736
rect -2990 748 -2984 1724
rect -2950 748 -2944 1724
rect -2990 736 -2944 748
rect -2732 1724 -2686 1736
rect -2732 748 -2726 1724
rect -2692 748 -2686 1724
rect -2732 736 -2686 748
rect -2474 1724 -2428 1736
rect -2474 748 -2468 1724
rect -2434 748 -2428 1724
rect -2474 736 -2428 748
rect -2216 1724 -2170 1736
rect -2216 748 -2210 1724
rect -2176 748 -2170 1724
rect -2216 736 -2170 748
rect -1958 1724 -1912 1736
rect -1958 748 -1952 1724
rect -1918 748 -1912 1724
rect -1958 736 -1912 748
rect -1700 1724 -1654 1736
rect -1700 748 -1694 1724
rect -1660 748 -1654 1724
rect -1700 736 -1654 748
rect -1442 1724 -1396 1736
rect -1442 748 -1436 1724
rect -1402 748 -1396 1724
rect -1442 736 -1396 748
rect -1184 1724 -1138 1736
rect -1184 748 -1178 1724
rect -1144 748 -1138 1724
rect -1184 736 -1138 748
rect -926 1724 -880 1736
rect -926 748 -920 1724
rect -886 748 -880 1724
rect -926 736 -880 748
rect -668 1724 -622 1736
rect -668 748 -662 1724
rect -628 748 -622 1724
rect -668 736 -622 748
rect -410 1724 -364 1736
rect -410 748 -404 1724
rect -370 748 -364 1724
rect -410 736 -364 748
rect -152 1724 -106 1736
rect -152 748 -146 1724
rect -112 748 -106 1724
rect -152 736 -106 748
rect 106 1724 152 1736
rect 106 748 112 1724
rect 146 748 152 1724
rect 106 736 152 748
rect 364 1724 410 1736
rect 364 748 370 1724
rect 404 748 410 1724
rect 364 736 410 748
rect 622 1724 668 1736
rect 622 748 628 1724
rect 662 748 668 1724
rect 622 736 668 748
rect 880 1724 926 1736
rect 880 748 886 1724
rect 920 748 926 1724
rect 880 736 926 748
rect 1138 1724 1184 1736
rect 1138 748 1144 1724
rect 1178 748 1184 1724
rect 1138 736 1184 748
rect 1396 1724 1442 1736
rect 1396 748 1402 1724
rect 1436 748 1442 1724
rect 1396 736 1442 748
rect 1654 1724 1700 1736
rect 1654 748 1660 1724
rect 1694 748 1700 1724
rect 1654 736 1700 748
rect 1912 1724 1958 1736
rect 1912 748 1918 1724
rect 1952 748 1958 1724
rect 1912 736 1958 748
rect 2170 1724 2216 1736
rect 2170 748 2176 1724
rect 2210 748 2216 1724
rect 2170 736 2216 748
rect 2428 1724 2474 1736
rect 2428 748 2434 1724
rect 2468 748 2474 1724
rect 2428 736 2474 748
rect 2686 1724 2732 1736
rect 2686 748 2692 1724
rect 2726 748 2732 1724
rect 2686 736 2732 748
rect 2944 1724 2990 1736
rect 2944 748 2950 1724
rect 2984 748 2990 1724
rect 2944 736 2990 748
rect -2934 689 -2742 695
rect -2934 655 -2922 689
rect -2754 655 -2742 689
rect -2934 649 -2742 655
rect -2676 689 -2484 695
rect -2676 655 -2664 689
rect -2496 655 -2484 689
rect -2676 649 -2484 655
rect -2418 689 -2226 695
rect -2418 655 -2406 689
rect -2238 655 -2226 689
rect -2418 649 -2226 655
rect -2160 689 -1968 695
rect -2160 655 -2148 689
rect -1980 655 -1968 689
rect -2160 649 -1968 655
rect -1902 689 -1710 695
rect -1902 655 -1890 689
rect -1722 655 -1710 689
rect -1902 649 -1710 655
rect -1644 689 -1452 695
rect -1644 655 -1632 689
rect -1464 655 -1452 689
rect -1644 649 -1452 655
rect -1386 689 -1194 695
rect -1386 655 -1374 689
rect -1206 655 -1194 689
rect -1386 649 -1194 655
rect -1128 689 -936 695
rect -1128 655 -1116 689
rect -948 655 -936 689
rect -1128 649 -936 655
rect -870 689 -678 695
rect -870 655 -858 689
rect -690 655 -678 689
rect -870 649 -678 655
rect -612 689 -420 695
rect -612 655 -600 689
rect -432 655 -420 689
rect -612 649 -420 655
rect -354 689 -162 695
rect -354 655 -342 689
rect -174 655 -162 689
rect -354 649 -162 655
rect -96 689 96 695
rect -96 655 -84 689
rect 84 655 96 689
rect -96 649 96 655
rect 162 689 354 695
rect 162 655 174 689
rect 342 655 354 689
rect 162 649 354 655
rect 420 689 612 695
rect 420 655 432 689
rect 600 655 612 689
rect 420 649 612 655
rect 678 689 870 695
rect 678 655 690 689
rect 858 655 870 689
rect 678 649 870 655
rect 936 689 1128 695
rect 936 655 948 689
rect 1116 655 1128 689
rect 936 649 1128 655
rect 1194 689 1386 695
rect 1194 655 1206 689
rect 1374 655 1386 689
rect 1194 649 1386 655
rect 1452 689 1644 695
rect 1452 655 1464 689
rect 1632 655 1644 689
rect 1452 649 1644 655
rect 1710 689 1902 695
rect 1710 655 1722 689
rect 1890 655 1902 689
rect 1710 649 1902 655
rect 1968 689 2160 695
rect 1968 655 1980 689
rect 2148 655 2160 689
rect 1968 649 2160 655
rect 2226 689 2418 695
rect 2226 655 2238 689
rect 2406 655 2418 689
rect 2226 649 2418 655
rect 2484 689 2676 695
rect 2484 655 2496 689
rect 2664 655 2676 689
rect 2484 649 2676 655
rect 2742 689 2934 695
rect 2742 655 2754 689
rect 2922 655 2934 689
rect 2742 649 2934 655
rect -2934 581 -2742 587
rect -2934 547 -2922 581
rect -2754 547 -2742 581
rect -2934 541 -2742 547
rect -2676 581 -2484 587
rect -2676 547 -2664 581
rect -2496 547 -2484 581
rect -2676 541 -2484 547
rect -2418 581 -2226 587
rect -2418 547 -2406 581
rect -2238 547 -2226 581
rect -2418 541 -2226 547
rect -2160 581 -1968 587
rect -2160 547 -2148 581
rect -1980 547 -1968 581
rect -2160 541 -1968 547
rect -1902 581 -1710 587
rect -1902 547 -1890 581
rect -1722 547 -1710 581
rect -1902 541 -1710 547
rect -1644 581 -1452 587
rect -1644 547 -1632 581
rect -1464 547 -1452 581
rect -1644 541 -1452 547
rect -1386 581 -1194 587
rect -1386 547 -1374 581
rect -1206 547 -1194 581
rect -1386 541 -1194 547
rect -1128 581 -936 587
rect -1128 547 -1116 581
rect -948 547 -936 581
rect -1128 541 -936 547
rect -870 581 -678 587
rect -870 547 -858 581
rect -690 547 -678 581
rect -870 541 -678 547
rect -612 581 -420 587
rect -612 547 -600 581
rect -432 547 -420 581
rect -612 541 -420 547
rect -354 581 -162 587
rect -354 547 -342 581
rect -174 547 -162 581
rect -354 541 -162 547
rect -96 581 96 587
rect -96 547 -84 581
rect 84 547 96 581
rect -96 541 96 547
rect 162 581 354 587
rect 162 547 174 581
rect 342 547 354 581
rect 162 541 354 547
rect 420 581 612 587
rect 420 547 432 581
rect 600 547 612 581
rect 420 541 612 547
rect 678 581 870 587
rect 678 547 690 581
rect 858 547 870 581
rect 678 541 870 547
rect 936 581 1128 587
rect 936 547 948 581
rect 1116 547 1128 581
rect 936 541 1128 547
rect 1194 581 1386 587
rect 1194 547 1206 581
rect 1374 547 1386 581
rect 1194 541 1386 547
rect 1452 581 1644 587
rect 1452 547 1464 581
rect 1632 547 1644 581
rect 1452 541 1644 547
rect 1710 581 1902 587
rect 1710 547 1722 581
rect 1890 547 1902 581
rect 1710 541 1902 547
rect 1968 581 2160 587
rect 1968 547 1980 581
rect 2148 547 2160 581
rect 1968 541 2160 547
rect 2226 581 2418 587
rect 2226 547 2238 581
rect 2406 547 2418 581
rect 2226 541 2418 547
rect 2484 581 2676 587
rect 2484 547 2496 581
rect 2664 547 2676 581
rect 2484 541 2676 547
rect 2742 581 2934 587
rect 2742 547 2754 581
rect 2922 547 2934 581
rect 2742 541 2934 547
rect -2990 488 -2944 500
rect -2990 -488 -2984 488
rect -2950 -488 -2944 488
rect -2990 -500 -2944 -488
rect -2732 488 -2686 500
rect -2732 -488 -2726 488
rect -2692 -488 -2686 488
rect -2732 -500 -2686 -488
rect -2474 488 -2428 500
rect -2474 -488 -2468 488
rect -2434 -488 -2428 488
rect -2474 -500 -2428 -488
rect -2216 488 -2170 500
rect -2216 -488 -2210 488
rect -2176 -488 -2170 488
rect -2216 -500 -2170 -488
rect -1958 488 -1912 500
rect -1958 -488 -1952 488
rect -1918 -488 -1912 488
rect -1958 -500 -1912 -488
rect -1700 488 -1654 500
rect -1700 -488 -1694 488
rect -1660 -488 -1654 488
rect -1700 -500 -1654 -488
rect -1442 488 -1396 500
rect -1442 -488 -1436 488
rect -1402 -488 -1396 488
rect -1442 -500 -1396 -488
rect -1184 488 -1138 500
rect -1184 -488 -1178 488
rect -1144 -488 -1138 488
rect -1184 -500 -1138 -488
rect -926 488 -880 500
rect -926 -488 -920 488
rect -886 -488 -880 488
rect -926 -500 -880 -488
rect -668 488 -622 500
rect -668 -488 -662 488
rect -628 -488 -622 488
rect -668 -500 -622 -488
rect -410 488 -364 500
rect -410 -488 -404 488
rect -370 -488 -364 488
rect -410 -500 -364 -488
rect -152 488 -106 500
rect -152 -488 -146 488
rect -112 -488 -106 488
rect -152 -500 -106 -488
rect 106 488 152 500
rect 106 -488 112 488
rect 146 -488 152 488
rect 106 -500 152 -488
rect 364 488 410 500
rect 364 -488 370 488
rect 404 -488 410 488
rect 364 -500 410 -488
rect 622 488 668 500
rect 622 -488 628 488
rect 662 -488 668 488
rect 622 -500 668 -488
rect 880 488 926 500
rect 880 -488 886 488
rect 920 -488 926 488
rect 880 -500 926 -488
rect 1138 488 1184 500
rect 1138 -488 1144 488
rect 1178 -488 1184 488
rect 1138 -500 1184 -488
rect 1396 488 1442 500
rect 1396 -488 1402 488
rect 1436 -488 1442 488
rect 1396 -500 1442 -488
rect 1654 488 1700 500
rect 1654 -488 1660 488
rect 1694 -488 1700 488
rect 1654 -500 1700 -488
rect 1912 488 1958 500
rect 1912 -488 1918 488
rect 1952 -488 1958 488
rect 1912 -500 1958 -488
rect 2170 488 2216 500
rect 2170 -488 2176 488
rect 2210 -488 2216 488
rect 2170 -500 2216 -488
rect 2428 488 2474 500
rect 2428 -488 2434 488
rect 2468 -488 2474 488
rect 2428 -500 2474 -488
rect 2686 488 2732 500
rect 2686 -488 2692 488
rect 2726 -488 2732 488
rect 2686 -500 2732 -488
rect 2944 488 2990 500
rect 2944 -488 2950 488
rect 2984 -488 2990 488
rect 2944 -500 2990 -488
rect -2934 -547 -2742 -541
rect -2934 -581 -2922 -547
rect -2754 -581 -2742 -547
rect -2934 -587 -2742 -581
rect -2676 -547 -2484 -541
rect -2676 -581 -2664 -547
rect -2496 -581 -2484 -547
rect -2676 -587 -2484 -581
rect -2418 -547 -2226 -541
rect -2418 -581 -2406 -547
rect -2238 -581 -2226 -547
rect -2418 -587 -2226 -581
rect -2160 -547 -1968 -541
rect -2160 -581 -2148 -547
rect -1980 -581 -1968 -547
rect -2160 -587 -1968 -581
rect -1902 -547 -1710 -541
rect -1902 -581 -1890 -547
rect -1722 -581 -1710 -547
rect -1902 -587 -1710 -581
rect -1644 -547 -1452 -541
rect -1644 -581 -1632 -547
rect -1464 -581 -1452 -547
rect -1644 -587 -1452 -581
rect -1386 -547 -1194 -541
rect -1386 -581 -1374 -547
rect -1206 -581 -1194 -547
rect -1386 -587 -1194 -581
rect -1128 -547 -936 -541
rect -1128 -581 -1116 -547
rect -948 -581 -936 -547
rect -1128 -587 -936 -581
rect -870 -547 -678 -541
rect -870 -581 -858 -547
rect -690 -581 -678 -547
rect -870 -587 -678 -581
rect -612 -547 -420 -541
rect -612 -581 -600 -547
rect -432 -581 -420 -547
rect -612 -587 -420 -581
rect -354 -547 -162 -541
rect -354 -581 -342 -547
rect -174 -581 -162 -547
rect -354 -587 -162 -581
rect -96 -547 96 -541
rect -96 -581 -84 -547
rect 84 -581 96 -547
rect -96 -587 96 -581
rect 162 -547 354 -541
rect 162 -581 174 -547
rect 342 -581 354 -547
rect 162 -587 354 -581
rect 420 -547 612 -541
rect 420 -581 432 -547
rect 600 -581 612 -547
rect 420 -587 612 -581
rect 678 -547 870 -541
rect 678 -581 690 -547
rect 858 -581 870 -547
rect 678 -587 870 -581
rect 936 -547 1128 -541
rect 936 -581 948 -547
rect 1116 -581 1128 -547
rect 936 -587 1128 -581
rect 1194 -547 1386 -541
rect 1194 -581 1206 -547
rect 1374 -581 1386 -547
rect 1194 -587 1386 -581
rect 1452 -547 1644 -541
rect 1452 -581 1464 -547
rect 1632 -581 1644 -547
rect 1452 -587 1644 -581
rect 1710 -547 1902 -541
rect 1710 -581 1722 -547
rect 1890 -581 1902 -547
rect 1710 -587 1902 -581
rect 1968 -547 2160 -541
rect 1968 -581 1980 -547
rect 2148 -581 2160 -547
rect 1968 -587 2160 -581
rect 2226 -547 2418 -541
rect 2226 -581 2238 -547
rect 2406 -581 2418 -547
rect 2226 -587 2418 -581
rect 2484 -547 2676 -541
rect 2484 -581 2496 -547
rect 2664 -581 2676 -547
rect 2484 -587 2676 -581
rect 2742 -547 2934 -541
rect 2742 -581 2754 -547
rect 2922 -581 2934 -547
rect 2742 -587 2934 -581
rect -2934 -655 -2742 -649
rect -2934 -689 -2922 -655
rect -2754 -689 -2742 -655
rect -2934 -695 -2742 -689
rect -2676 -655 -2484 -649
rect -2676 -689 -2664 -655
rect -2496 -689 -2484 -655
rect -2676 -695 -2484 -689
rect -2418 -655 -2226 -649
rect -2418 -689 -2406 -655
rect -2238 -689 -2226 -655
rect -2418 -695 -2226 -689
rect -2160 -655 -1968 -649
rect -2160 -689 -2148 -655
rect -1980 -689 -1968 -655
rect -2160 -695 -1968 -689
rect -1902 -655 -1710 -649
rect -1902 -689 -1890 -655
rect -1722 -689 -1710 -655
rect -1902 -695 -1710 -689
rect -1644 -655 -1452 -649
rect -1644 -689 -1632 -655
rect -1464 -689 -1452 -655
rect -1644 -695 -1452 -689
rect -1386 -655 -1194 -649
rect -1386 -689 -1374 -655
rect -1206 -689 -1194 -655
rect -1386 -695 -1194 -689
rect -1128 -655 -936 -649
rect -1128 -689 -1116 -655
rect -948 -689 -936 -655
rect -1128 -695 -936 -689
rect -870 -655 -678 -649
rect -870 -689 -858 -655
rect -690 -689 -678 -655
rect -870 -695 -678 -689
rect -612 -655 -420 -649
rect -612 -689 -600 -655
rect -432 -689 -420 -655
rect -612 -695 -420 -689
rect -354 -655 -162 -649
rect -354 -689 -342 -655
rect -174 -689 -162 -655
rect -354 -695 -162 -689
rect -96 -655 96 -649
rect -96 -689 -84 -655
rect 84 -689 96 -655
rect -96 -695 96 -689
rect 162 -655 354 -649
rect 162 -689 174 -655
rect 342 -689 354 -655
rect 162 -695 354 -689
rect 420 -655 612 -649
rect 420 -689 432 -655
rect 600 -689 612 -655
rect 420 -695 612 -689
rect 678 -655 870 -649
rect 678 -689 690 -655
rect 858 -689 870 -655
rect 678 -695 870 -689
rect 936 -655 1128 -649
rect 936 -689 948 -655
rect 1116 -689 1128 -655
rect 936 -695 1128 -689
rect 1194 -655 1386 -649
rect 1194 -689 1206 -655
rect 1374 -689 1386 -655
rect 1194 -695 1386 -689
rect 1452 -655 1644 -649
rect 1452 -689 1464 -655
rect 1632 -689 1644 -655
rect 1452 -695 1644 -689
rect 1710 -655 1902 -649
rect 1710 -689 1722 -655
rect 1890 -689 1902 -655
rect 1710 -695 1902 -689
rect 1968 -655 2160 -649
rect 1968 -689 1980 -655
rect 2148 -689 2160 -655
rect 1968 -695 2160 -689
rect 2226 -655 2418 -649
rect 2226 -689 2238 -655
rect 2406 -689 2418 -655
rect 2226 -695 2418 -689
rect 2484 -655 2676 -649
rect 2484 -689 2496 -655
rect 2664 -689 2676 -655
rect 2484 -695 2676 -689
rect 2742 -655 2934 -649
rect 2742 -689 2754 -655
rect 2922 -689 2934 -655
rect 2742 -695 2934 -689
rect -2990 -748 -2944 -736
rect -2990 -1724 -2984 -748
rect -2950 -1724 -2944 -748
rect -2990 -1736 -2944 -1724
rect -2732 -748 -2686 -736
rect -2732 -1724 -2726 -748
rect -2692 -1724 -2686 -748
rect -2732 -1736 -2686 -1724
rect -2474 -748 -2428 -736
rect -2474 -1724 -2468 -748
rect -2434 -1724 -2428 -748
rect -2474 -1736 -2428 -1724
rect -2216 -748 -2170 -736
rect -2216 -1724 -2210 -748
rect -2176 -1724 -2170 -748
rect -2216 -1736 -2170 -1724
rect -1958 -748 -1912 -736
rect -1958 -1724 -1952 -748
rect -1918 -1724 -1912 -748
rect -1958 -1736 -1912 -1724
rect -1700 -748 -1654 -736
rect -1700 -1724 -1694 -748
rect -1660 -1724 -1654 -748
rect -1700 -1736 -1654 -1724
rect -1442 -748 -1396 -736
rect -1442 -1724 -1436 -748
rect -1402 -1724 -1396 -748
rect -1442 -1736 -1396 -1724
rect -1184 -748 -1138 -736
rect -1184 -1724 -1178 -748
rect -1144 -1724 -1138 -748
rect -1184 -1736 -1138 -1724
rect -926 -748 -880 -736
rect -926 -1724 -920 -748
rect -886 -1724 -880 -748
rect -926 -1736 -880 -1724
rect -668 -748 -622 -736
rect -668 -1724 -662 -748
rect -628 -1724 -622 -748
rect -668 -1736 -622 -1724
rect -410 -748 -364 -736
rect -410 -1724 -404 -748
rect -370 -1724 -364 -748
rect -410 -1736 -364 -1724
rect -152 -748 -106 -736
rect -152 -1724 -146 -748
rect -112 -1724 -106 -748
rect -152 -1736 -106 -1724
rect 106 -748 152 -736
rect 106 -1724 112 -748
rect 146 -1724 152 -748
rect 106 -1736 152 -1724
rect 364 -748 410 -736
rect 364 -1724 370 -748
rect 404 -1724 410 -748
rect 364 -1736 410 -1724
rect 622 -748 668 -736
rect 622 -1724 628 -748
rect 662 -1724 668 -748
rect 622 -1736 668 -1724
rect 880 -748 926 -736
rect 880 -1724 886 -748
rect 920 -1724 926 -748
rect 880 -1736 926 -1724
rect 1138 -748 1184 -736
rect 1138 -1724 1144 -748
rect 1178 -1724 1184 -748
rect 1138 -1736 1184 -1724
rect 1396 -748 1442 -736
rect 1396 -1724 1402 -748
rect 1436 -1724 1442 -748
rect 1396 -1736 1442 -1724
rect 1654 -748 1700 -736
rect 1654 -1724 1660 -748
rect 1694 -1724 1700 -748
rect 1654 -1736 1700 -1724
rect 1912 -748 1958 -736
rect 1912 -1724 1918 -748
rect 1952 -1724 1958 -748
rect 1912 -1736 1958 -1724
rect 2170 -748 2216 -736
rect 2170 -1724 2176 -748
rect 2210 -1724 2216 -748
rect 2170 -1736 2216 -1724
rect 2428 -748 2474 -736
rect 2428 -1724 2434 -748
rect 2468 -1724 2474 -748
rect 2428 -1736 2474 -1724
rect 2686 -748 2732 -736
rect 2686 -1724 2692 -748
rect 2726 -1724 2732 -748
rect 2686 -1736 2732 -1724
rect 2944 -748 2990 -736
rect 2944 -1724 2950 -748
rect 2984 -1724 2990 -748
rect 2944 -1736 2990 -1724
rect -2934 -1783 -2742 -1777
rect -2934 -1817 -2922 -1783
rect -2754 -1817 -2742 -1783
rect -2934 -1823 -2742 -1817
rect -2676 -1783 -2484 -1777
rect -2676 -1817 -2664 -1783
rect -2496 -1817 -2484 -1783
rect -2676 -1823 -2484 -1817
rect -2418 -1783 -2226 -1777
rect -2418 -1817 -2406 -1783
rect -2238 -1817 -2226 -1783
rect -2418 -1823 -2226 -1817
rect -2160 -1783 -1968 -1777
rect -2160 -1817 -2148 -1783
rect -1980 -1817 -1968 -1783
rect -2160 -1823 -1968 -1817
rect -1902 -1783 -1710 -1777
rect -1902 -1817 -1890 -1783
rect -1722 -1817 -1710 -1783
rect -1902 -1823 -1710 -1817
rect -1644 -1783 -1452 -1777
rect -1644 -1817 -1632 -1783
rect -1464 -1817 -1452 -1783
rect -1644 -1823 -1452 -1817
rect -1386 -1783 -1194 -1777
rect -1386 -1817 -1374 -1783
rect -1206 -1817 -1194 -1783
rect -1386 -1823 -1194 -1817
rect -1128 -1783 -936 -1777
rect -1128 -1817 -1116 -1783
rect -948 -1817 -936 -1783
rect -1128 -1823 -936 -1817
rect -870 -1783 -678 -1777
rect -870 -1817 -858 -1783
rect -690 -1817 -678 -1783
rect -870 -1823 -678 -1817
rect -612 -1783 -420 -1777
rect -612 -1817 -600 -1783
rect -432 -1817 -420 -1783
rect -612 -1823 -420 -1817
rect -354 -1783 -162 -1777
rect -354 -1817 -342 -1783
rect -174 -1817 -162 -1783
rect -354 -1823 -162 -1817
rect -96 -1783 96 -1777
rect -96 -1817 -84 -1783
rect 84 -1817 96 -1783
rect -96 -1823 96 -1817
rect 162 -1783 354 -1777
rect 162 -1817 174 -1783
rect 342 -1817 354 -1783
rect 162 -1823 354 -1817
rect 420 -1783 612 -1777
rect 420 -1817 432 -1783
rect 600 -1817 612 -1783
rect 420 -1823 612 -1817
rect 678 -1783 870 -1777
rect 678 -1817 690 -1783
rect 858 -1817 870 -1783
rect 678 -1823 870 -1817
rect 936 -1783 1128 -1777
rect 936 -1817 948 -1783
rect 1116 -1817 1128 -1783
rect 936 -1823 1128 -1817
rect 1194 -1783 1386 -1777
rect 1194 -1817 1206 -1783
rect 1374 -1817 1386 -1783
rect 1194 -1823 1386 -1817
rect 1452 -1783 1644 -1777
rect 1452 -1817 1464 -1783
rect 1632 -1817 1644 -1783
rect 1452 -1823 1644 -1817
rect 1710 -1783 1902 -1777
rect 1710 -1817 1722 -1783
rect 1890 -1817 1902 -1783
rect 1710 -1823 1902 -1817
rect 1968 -1783 2160 -1777
rect 1968 -1817 1980 -1783
rect 2148 -1817 2160 -1783
rect 1968 -1823 2160 -1817
rect 2226 -1783 2418 -1777
rect 2226 -1817 2238 -1783
rect 2406 -1817 2418 -1783
rect 2226 -1823 2418 -1817
rect 2484 -1783 2676 -1777
rect 2484 -1817 2496 -1783
rect 2664 -1817 2676 -1783
rect 2484 -1823 2676 -1817
rect 2742 -1783 2934 -1777
rect 2742 -1817 2754 -1783
rect 2922 -1817 2934 -1783
rect 2742 -1823 2934 -1817
rect -2934 -1891 -2742 -1885
rect -2934 -1925 -2922 -1891
rect -2754 -1925 -2742 -1891
rect -2934 -1931 -2742 -1925
rect -2676 -1891 -2484 -1885
rect -2676 -1925 -2664 -1891
rect -2496 -1925 -2484 -1891
rect -2676 -1931 -2484 -1925
rect -2418 -1891 -2226 -1885
rect -2418 -1925 -2406 -1891
rect -2238 -1925 -2226 -1891
rect -2418 -1931 -2226 -1925
rect -2160 -1891 -1968 -1885
rect -2160 -1925 -2148 -1891
rect -1980 -1925 -1968 -1891
rect -2160 -1931 -1968 -1925
rect -1902 -1891 -1710 -1885
rect -1902 -1925 -1890 -1891
rect -1722 -1925 -1710 -1891
rect -1902 -1931 -1710 -1925
rect -1644 -1891 -1452 -1885
rect -1644 -1925 -1632 -1891
rect -1464 -1925 -1452 -1891
rect -1644 -1931 -1452 -1925
rect -1386 -1891 -1194 -1885
rect -1386 -1925 -1374 -1891
rect -1206 -1925 -1194 -1891
rect -1386 -1931 -1194 -1925
rect -1128 -1891 -936 -1885
rect -1128 -1925 -1116 -1891
rect -948 -1925 -936 -1891
rect -1128 -1931 -936 -1925
rect -870 -1891 -678 -1885
rect -870 -1925 -858 -1891
rect -690 -1925 -678 -1891
rect -870 -1931 -678 -1925
rect -612 -1891 -420 -1885
rect -612 -1925 -600 -1891
rect -432 -1925 -420 -1891
rect -612 -1931 -420 -1925
rect -354 -1891 -162 -1885
rect -354 -1925 -342 -1891
rect -174 -1925 -162 -1891
rect -354 -1931 -162 -1925
rect -96 -1891 96 -1885
rect -96 -1925 -84 -1891
rect 84 -1925 96 -1891
rect -96 -1931 96 -1925
rect 162 -1891 354 -1885
rect 162 -1925 174 -1891
rect 342 -1925 354 -1891
rect 162 -1931 354 -1925
rect 420 -1891 612 -1885
rect 420 -1925 432 -1891
rect 600 -1925 612 -1891
rect 420 -1931 612 -1925
rect 678 -1891 870 -1885
rect 678 -1925 690 -1891
rect 858 -1925 870 -1891
rect 678 -1931 870 -1925
rect 936 -1891 1128 -1885
rect 936 -1925 948 -1891
rect 1116 -1925 1128 -1891
rect 936 -1931 1128 -1925
rect 1194 -1891 1386 -1885
rect 1194 -1925 1206 -1891
rect 1374 -1925 1386 -1891
rect 1194 -1931 1386 -1925
rect 1452 -1891 1644 -1885
rect 1452 -1925 1464 -1891
rect 1632 -1925 1644 -1891
rect 1452 -1931 1644 -1925
rect 1710 -1891 1902 -1885
rect 1710 -1925 1722 -1891
rect 1890 -1925 1902 -1891
rect 1710 -1931 1902 -1925
rect 1968 -1891 2160 -1885
rect 1968 -1925 1980 -1891
rect 2148 -1925 2160 -1891
rect 1968 -1931 2160 -1925
rect 2226 -1891 2418 -1885
rect 2226 -1925 2238 -1891
rect 2406 -1925 2418 -1891
rect 2226 -1931 2418 -1925
rect 2484 -1891 2676 -1885
rect 2484 -1925 2496 -1891
rect 2664 -1925 2676 -1891
rect 2484 -1931 2676 -1925
rect 2742 -1891 2934 -1885
rect 2742 -1925 2754 -1891
rect 2922 -1925 2934 -1891
rect 2742 -1931 2934 -1925
rect -2990 -1984 -2944 -1972
rect -2990 -2960 -2984 -1984
rect -2950 -2960 -2944 -1984
rect -2990 -2972 -2944 -2960
rect -2732 -1984 -2686 -1972
rect -2732 -2960 -2726 -1984
rect -2692 -2960 -2686 -1984
rect -2732 -2972 -2686 -2960
rect -2474 -1984 -2428 -1972
rect -2474 -2960 -2468 -1984
rect -2434 -2960 -2428 -1984
rect -2474 -2972 -2428 -2960
rect -2216 -1984 -2170 -1972
rect -2216 -2960 -2210 -1984
rect -2176 -2960 -2170 -1984
rect -2216 -2972 -2170 -2960
rect -1958 -1984 -1912 -1972
rect -1958 -2960 -1952 -1984
rect -1918 -2960 -1912 -1984
rect -1958 -2972 -1912 -2960
rect -1700 -1984 -1654 -1972
rect -1700 -2960 -1694 -1984
rect -1660 -2960 -1654 -1984
rect -1700 -2972 -1654 -2960
rect -1442 -1984 -1396 -1972
rect -1442 -2960 -1436 -1984
rect -1402 -2960 -1396 -1984
rect -1442 -2972 -1396 -2960
rect -1184 -1984 -1138 -1972
rect -1184 -2960 -1178 -1984
rect -1144 -2960 -1138 -1984
rect -1184 -2972 -1138 -2960
rect -926 -1984 -880 -1972
rect -926 -2960 -920 -1984
rect -886 -2960 -880 -1984
rect -926 -2972 -880 -2960
rect -668 -1984 -622 -1972
rect -668 -2960 -662 -1984
rect -628 -2960 -622 -1984
rect -668 -2972 -622 -2960
rect -410 -1984 -364 -1972
rect -410 -2960 -404 -1984
rect -370 -2960 -364 -1984
rect -410 -2972 -364 -2960
rect -152 -1984 -106 -1972
rect -152 -2960 -146 -1984
rect -112 -2960 -106 -1984
rect -152 -2972 -106 -2960
rect 106 -1984 152 -1972
rect 106 -2960 112 -1984
rect 146 -2960 152 -1984
rect 106 -2972 152 -2960
rect 364 -1984 410 -1972
rect 364 -2960 370 -1984
rect 404 -2960 410 -1984
rect 364 -2972 410 -2960
rect 622 -1984 668 -1972
rect 622 -2960 628 -1984
rect 662 -2960 668 -1984
rect 622 -2972 668 -2960
rect 880 -1984 926 -1972
rect 880 -2960 886 -1984
rect 920 -2960 926 -1984
rect 880 -2972 926 -2960
rect 1138 -1984 1184 -1972
rect 1138 -2960 1144 -1984
rect 1178 -2960 1184 -1984
rect 1138 -2972 1184 -2960
rect 1396 -1984 1442 -1972
rect 1396 -2960 1402 -1984
rect 1436 -2960 1442 -1984
rect 1396 -2972 1442 -2960
rect 1654 -1984 1700 -1972
rect 1654 -2960 1660 -1984
rect 1694 -2960 1700 -1984
rect 1654 -2972 1700 -2960
rect 1912 -1984 1958 -1972
rect 1912 -2960 1918 -1984
rect 1952 -2960 1958 -1984
rect 1912 -2972 1958 -2960
rect 2170 -1984 2216 -1972
rect 2170 -2960 2176 -1984
rect 2210 -2960 2216 -1984
rect 2170 -2972 2216 -2960
rect 2428 -1984 2474 -1972
rect 2428 -2960 2434 -1984
rect 2468 -2960 2474 -1984
rect 2428 -2972 2474 -2960
rect 2686 -1984 2732 -1972
rect 2686 -2960 2692 -1984
rect 2726 -2960 2732 -1984
rect 2686 -2972 2732 -2960
rect 2944 -1984 2990 -1972
rect 2944 -2960 2950 -1984
rect 2984 -2960 2990 -1984
rect 2944 -2972 2990 -2960
rect -2934 -3019 -2742 -3013
rect -2934 -3053 -2922 -3019
rect -2754 -3053 -2742 -3019
rect -2934 -3059 -2742 -3053
rect -2676 -3019 -2484 -3013
rect -2676 -3053 -2664 -3019
rect -2496 -3053 -2484 -3019
rect -2676 -3059 -2484 -3053
rect -2418 -3019 -2226 -3013
rect -2418 -3053 -2406 -3019
rect -2238 -3053 -2226 -3019
rect -2418 -3059 -2226 -3053
rect -2160 -3019 -1968 -3013
rect -2160 -3053 -2148 -3019
rect -1980 -3053 -1968 -3019
rect -2160 -3059 -1968 -3053
rect -1902 -3019 -1710 -3013
rect -1902 -3053 -1890 -3019
rect -1722 -3053 -1710 -3019
rect -1902 -3059 -1710 -3053
rect -1644 -3019 -1452 -3013
rect -1644 -3053 -1632 -3019
rect -1464 -3053 -1452 -3019
rect -1644 -3059 -1452 -3053
rect -1386 -3019 -1194 -3013
rect -1386 -3053 -1374 -3019
rect -1206 -3053 -1194 -3019
rect -1386 -3059 -1194 -3053
rect -1128 -3019 -936 -3013
rect -1128 -3053 -1116 -3019
rect -948 -3053 -936 -3019
rect -1128 -3059 -936 -3053
rect -870 -3019 -678 -3013
rect -870 -3053 -858 -3019
rect -690 -3053 -678 -3019
rect -870 -3059 -678 -3053
rect -612 -3019 -420 -3013
rect -612 -3053 -600 -3019
rect -432 -3053 -420 -3019
rect -612 -3059 -420 -3053
rect -354 -3019 -162 -3013
rect -354 -3053 -342 -3019
rect -174 -3053 -162 -3019
rect -354 -3059 -162 -3053
rect -96 -3019 96 -3013
rect -96 -3053 -84 -3019
rect 84 -3053 96 -3019
rect -96 -3059 96 -3053
rect 162 -3019 354 -3013
rect 162 -3053 174 -3019
rect 342 -3053 354 -3019
rect 162 -3059 354 -3053
rect 420 -3019 612 -3013
rect 420 -3053 432 -3019
rect 600 -3053 612 -3019
rect 420 -3059 612 -3053
rect 678 -3019 870 -3013
rect 678 -3053 690 -3019
rect 858 -3053 870 -3019
rect 678 -3059 870 -3053
rect 936 -3019 1128 -3013
rect 936 -3053 948 -3019
rect 1116 -3053 1128 -3019
rect 936 -3059 1128 -3053
rect 1194 -3019 1386 -3013
rect 1194 -3053 1206 -3019
rect 1374 -3053 1386 -3019
rect 1194 -3059 1386 -3053
rect 1452 -3019 1644 -3013
rect 1452 -3053 1464 -3019
rect 1632 -3053 1644 -3019
rect 1452 -3059 1644 -3053
rect 1710 -3019 1902 -3013
rect 1710 -3053 1722 -3019
rect 1890 -3053 1902 -3019
rect 1710 -3059 1902 -3053
rect 1968 -3019 2160 -3013
rect 1968 -3053 1980 -3019
rect 2148 -3053 2160 -3019
rect 1968 -3059 2160 -3053
rect 2226 -3019 2418 -3013
rect 2226 -3053 2238 -3019
rect 2406 -3053 2418 -3019
rect 2226 -3059 2418 -3053
rect 2484 -3019 2676 -3013
rect 2484 -3053 2496 -3019
rect 2664 -3053 2676 -3019
rect 2484 -3059 2676 -3053
rect 2742 -3019 2934 -3013
rect 2742 -3053 2754 -3019
rect 2922 -3053 2934 -3019
rect 2742 -3059 2934 -3053
<< properties >>
string FIXED_BBOX -3101 -3174 3101 3174
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 1 m 5 nf 23 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
